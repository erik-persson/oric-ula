//----------------------------------------------------------------------------
// Top - Extracted by tractor
//----------------------------------------------------------------------------

module Top
(
  input  wire    CLK,
  input  wire    A8,
  input  wire    A9,
  input  wire    A10,
  input  wire    A11,
  input  wire    A12,
  input  wire    A13,
  input  wire    A14,
  input  wire    A15,
  input  wire    D0,
  input  wire    D1,
  input  wire    D2,
  input  wire    D3,
  input  wire    D4,
  input  wire    D5,
  input  wire    D6,
  input  wire    D7,
  input  wire    RnW,
  input  wire    nMAP,
  output wire    RC0,
  output wire    RC1,
  output wire    RC2,
  output wire    RC3,
  output wire    RC4,
  output wire    RC5,
  output wire    RC6,
  output wire    RC7,
  output wire    MXSEL,
  output wire    nROM,
  output wire    PHI,
  output wire    CAS,
  output wire    RAS,
  output wire    WE,
  output wire    nIO,
  output wire    SYNC,
  output wire    RED,
  output wire    GREEN,
  output wire    BLUE
);

  wire    I_1039_D;
  wire    I_1089_D;
  wire    I_1091_D;
  reg     I_1093_D = 1'b1;
  reg     I_1095_D = 1'b1;
  wire    I_1103_D;
  wire    I_1111_D;
  wire    I_1115_D;
  reg     I_1119_D = 1'b1;
  wire    I_1185_D;
  wire    I_1211_D;
  wire    I_1213_D;
  wire    I_1251_D;
  reg     I_1253_D = 1'b1;
  reg     I_1255_D = 1'b1;
  reg     I_1257_D = 1'b1;
  reg     I_1259_D = 1'b1;
  wire    I_1265_D;
  reg     I_1267_D = 1'b1;
  reg     I_1269_D = 1'b1;
  reg     I_1271_D = 1'b1;
  wire    I_1275_D;
  wire    I_1279_D;
  wire    I_128_D;
  reg     I_133_D = 1'b1;
  wire    I_1359_D;
  reg     I_135_D = 1'b1;
  reg     I_1413_D = 1'b1;
  reg     I_1415_D = 1'b1;
  reg     I_1417_D = 1'b1;
  reg     I_1419_D = 1'b1;
  wire    I_1423_D;
  wire    I_1425_S;
  reg     I_1427_D = 1'b1;
  reg     I_1429_D = 1'b1;
  reg     I_1431_D = 1'b1;
  wire    I_1433_D;
  wire    I_1435_D;
  reg     I_1439_D = 1'b1;
  wire    I_1439_S;
  wire    I_1499_D;
  wire    I_1518_D;
  wire    I_1535_D;
  reg     I_153_D = 1'b1;
  wire    I_155_D;
  reg     I_1569_D = 1'b1;
  reg     I_1571_D = 1'b1;
  reg     I_1573_D = 1'b1;
  reg     I_1575_D = 1'b1;
  reg     I_157_D = 1'b1;
  wire    I_1585_D;
  reg     I_1591_D = 1'b1;
  reg     I_1593_D = 1'b1;
  wire    I_1648_D;
  wire    I_1673_D;
  wire    I_1679_D;
  wire    I_1693_D;
  wire    I_1695_D;
  reg     I_1729_D = 1'b1;
  reg     I_1731_D = 1'b1;
  reg     I_1733_D = 1'b1;
  reg     I_1735_D = 1'b1;
  wire    I_1737_D;
  wire    I_1743_D;
  wire    I_1807_D;
  wire    I_1832_D;
  wire    I_1845_D;
  wire    I_1855_D;
  wire    I_1889_D;
  wire    I_1891_S;
  reg     I_1893_D = 1'b1;
  reg     I_1895_D = 1'b1;
  wire    I_1899_S;
  wire    I_1901_D;
  reg     I_1911_D = 1'b1;
  reg     I_1913_D = 1'b1;
  wire    I_1913_S;
  wire    I_1915_S;
  wire    I_1917_D;
  wire    I_1962_D;
  wire    I_1987_D;
  wire    I_1999_D;
  wire    I_2011_D;
  wire    I_2013_D;
  wire    I_2015_D;
  reg     I_2049_D = 1'b1;
  wire    I_2051_D;
  reg     I_2053_D = 1'b1;
  reg     I_2055_D = 1'b1;
  wire    I_2063_D;
  wire    I_2065_S;
  wire    I_2069_D;
  wire    I_2071_D;
  wire    I_2071_S;
  reg     I_2073_D = 1'b1;
  wire    I_2075_D;
  wire    I_2077_D;
  wire    I_2115_D;
  wire    I_2127_D;
  wire    I_2132_D;
  wire    I_2139_D;
  wire    I_2154_D;
  wire    I_2173_D;
  wire    I_2175_D;
  reg     I_2209_D = 1'b1;
  wire    I_2211_D;
  reg     I_2213_D = 1'b1;
  reg     I_2215_D = 1'b1;
  wire    I_2225_D;
  wire    I_2231_S;
  reg     I_2233_D = 1'b1;
  wire    I_2235_D;
  wire    I_2237_D;
  wire    I_225_D;
  wire    I_2275_D;
  wire    I_227_D;
  wire    I_2288_D;
  wire    I_2319_D;
  wire    I_2331_D;
  wire    I_2333_D;
  wire    I_2335_D;
  wire    I_235_D;
  reg     I_2369_D = 1'b1;
  wire    I_2371_S;
  reg     I_2373_D = 1'b1;
  reg     I_2375_D = 1'b1;
  wire    I_2379_S;
  wire    I_2383_D;
  wire    I_2391_D;
  reg     I_2393_D = 1'b1;
  wire    I_2395_D;
  wire    I_2397_D;
  wire    I_2447_D;
  wire    I_2454_D;
  wire    I_2491_D;
  wire    I_2493_D;
  wire    I_2495_D;
  reg     I_2529_D = 1'b1;
  reg     I_2533_D = 1'b1;
  reg     I_2535_D = 1'b1;
  wire    I_2539_S;
  wire    I_2545_S;
  wire    I_2549_D;
  wire    I_2549_S;
  reg     I_2553_D = 1'b1;
  wire    I_2555_D;
  wire    I_2557_D;
  wire    I_2632_D;
  wire    I_2634_D;
  wire    I_2650_D;
  wire    I_2653_D;
  wire    I_2655_D;
  reg     I_2689_D = 1'b1;
  reg     I_2693_D = 1'b1;
  reg     I_2695_D = 1'b1;
  wire    I_2699_D;
  wire    I_2705_S;
  wire    I_2709_D;
  wire    I_2709_S;
  wire    I_2711_S;
  reg     I_2713_D = 1'b1;
  wire    I_2715_D;
  wire    I_2717_D;
  wire    I_2794_D;
  wire    I_2811_D;
  wire    I_2813_D;
  wire    I_2815_D;
  reg     I_2849_D = 1'b1;
  reg     I_2853_D = 1'b1;
  reg     I_2855_D = 1'b1;
  wire    I_2865_D;
  wire    I_2869_D;
  wire    I_2871_D;
  wire    I_2871_S;
  reg     I_2873_D = 1'b1;
  wire    I_2875_D;
  wire    I_2877_D;
  wire    I_289_D;
  wire    I_291_D;
  wire    I_2928_D;
  reg     I_293_D = 1'b1;
  wire    I_2953_D;
  wire    I_2955_D;
  wire    I_2957_D;
  reg     I_295_D = 1'b1;
  wire    I_2971_D;
  wire    I_2972_D;
  wire    I_2975_D;
  reg     I_3009_D = 1'b1;
  reg     I_3013_D = 1'b1;
  reg     I_3015_D = 1'b1;
  wire    I_3017_D;
  wire    I_3021_D;
  wire    I_3023_D;
  wire    I_3027_D;
  wire    I_3029_D;
  wire    I_3031_D;
  wire    I_3031_S;
  reg     I_3033_D = 1'b1;
  wire    I_3035_D;
  wire    I_3075_D;
  wire    I_3083_D;
  wire    I_3086_D;
  wire    I_3112_D;
  wire    I_3116_D;
  reg     I_311_D = 1'b1;
  wire    I_3130_D;
  wire    I_3133_D;
  wire    I_3135_D;
  reg     I_313_D = 1'b1;
  reg     I_3169_D = 1'b1;
  wire    I_3171_D;
  reg     I_3173_D = 1'b1;
  reg     I_3175_D = 1'b1;
  wire    I_3177_D;
  reg     I_317_D = 1'b1;
  wire    I_3185_S;
  wire    I_3189_S;
  wire    I_3191_D;
  wire    I_3191_S;
  wire    I_3193_D;
  wire    I_3197_D;
  reg     I_319_D = 1'b1;
  wire    I_3285_D;
  wire    I_3287_D;
  wire    I_3289_D;
  wire    I_3291_D;
  wire    I_3293_D;
  reg     I_3329_D = 1'b1;
  reg     I_3333_D = 1'b1;
  reg     I_3335_D = 1'b1;
  wire    I_3337_D;
  wire    I_3339_D;
  wire    I_3345_D;
  wire    I_3345_S;
  wire    I_3347_D;
  wire    I_3349_D;
  wire    I_3353_D;
  wire    I_3357_D;
  wire    I_3413_D;
  wire    I_3427_D;
  wire    I_3447_D;
  wire    I_3449_D;
  wire    I_3451_D;
  wire    I_3453_D;
  reg     I_3489_D = 1'b1;
  wire    I_3491_S;
  reg     I_3493_D = 1'b1;
  reg     I_3495_D = 1'b1;
  wire    I_3497_S;
  wire    I_3499_D;
  wire    I_3499_S;
  wire    I_3501_D;
  wire    I_3503_D;
  wire    I_3503_S;
  wire    I_3505_D;
  wire    I_3507_D;
  wire    I_3517_D;
  wire    I_355_D;
  wire    I_3562_D;
  wire    I_3565_D;
  wire    I_3568_D;
  wire    I_3585_D;
  wire    I_3587_D;
  wire    I_3607_D;
  wire    I_3609_D;
  wire    I_3611_D;
  wire    I_3613_D;
  wire    I_3615_D;
  reg     I_3653_D = 1'b1;
  reg     I_3655_D = 1'b1;
  wire    I_3663_D;
  wire    I_3663_S;
  wire    I_3667_D;
  wire    I_3669_D;
  wire    I_3669_S;
  wire    I_3677_D;
  wire    I_3725_D;
  wire    I_3745_D;
  wire    I_3747_D;
  wire    I_3753_D;
  wire    I_3755_S;
  wire    I_3767_D;
  wire    I_3769_D;
  wire    I_3771_D;
  wire    I_3773_D;
  wire    I_3775_D;
  wire    I_3809_D;
  wire    I_3811_D;
  reg     I_3813_D = 1'b1;
  reg     I_3815_D = 1'b1;
  wire    I_3817_D;
  wire    I_3823_D;
  wire    I_3823_S;
  wire    I_3825_D;
  wire    I_3825_S;
  wire    I_3827_D;
  wire    I_3829_D;
  wire    I_3829_S;
  wire    I_3831_D;
  wire    I_3835_D;
  wire    I_3837_D;
  wire    I_3883_D;
  wire    I_3884_D;
  wire    I_3904_D;
  wire    I_3906_D;
  wire    I_3909_D;
  wire    I_3911_D;
  wire    I_3913_S;
  wire    I_3926_D;
  wire    I_3929_D;
  wire    I_3931_D;
  wire    I_3933_D;
  wire    I_3935_D;
  wire    I_395_D;
  wire    I_3973_D;
  wire    I_3975_D;
  wire    I_3977_D;
  wire    I_3981_D;
  wire    I_3985_D;
  wire    I_3985_S;
  wire    I_3995_D;
  wire    I_3997_D;
  wire    I_448_D;
  reg     I_453_D = 1'b1;
  reg     I_455_D = 1'b1;
  wire    I_457_D;
  reg     I_471_D = 1'b1;
  reg     I_473_D = 1'b1;
  wire    I_475_D;
  wire    I_477_D;
  reg     I_479_D = 1'b1;
  wire    I_524_D;
  wire    I_545_D;
  wire    I_547_D;
  wire    I_553_D;
  wire    I_555_D;
  wire    I_573_D;
  wire    I_609_D;
  wire    I_611_D;
  reg     I_613_D = 1'b1;
  reg     I_615_D = 1'b1;
  wire    I_631_D;
  reg     I_633_D = 1'b1;
  reg     I_637_D = 1'b1;
  wire    I_675_D;
  wire    I_67_S;
  wire    I_715_D;
  wire    I_768_D;
  reg     I_773_D = 1'b1;
  reg     I_775_D = 1'b1;
  reg     I_777_D = 1'b1;
  reg     I_791_D = 1'b1;
  reg     I_793_D = 1'b1;
  wire    I_795_D;
  reg     I_797_D = 1'b1;
  wire    I_865_D;
  wire    I_867_D;
  wire    I_929_D;
  wire    I_931_D;
  reg     I_933_D = 1'b1;
  reg     I_935_D = 1'b1;
  reg     I_937_D = 1'b1;
  reg     I_951_D = 1'b1;
  reg     I_953_D = 1'b1;
  wire    I_957_D;
  reg     I_959_D = 1'b1;
  wire    I_995_D;

  assign RC0 = I_3677_D;
  assign RC1 = I_3995_D;
  assign RC2 = I_3353_D;
  assign RC3 = I_2077_D;
  assign RC4 = I_2397_D;
  assign RC5 = I_2717_D;
  assign RC6 = I_2972_D;
  assign RC7 = I_3357_D;
  assign MXSEL = I_1915_S;
  assign nROM = I_3884_D;
  assign PHI = !I_1119_D;
  assign CAS = !I_1115_D;
  assign RAS = I_1427_D;
  assign WE = !I_3981_D;
  assign nIO = !I_3755_S;
  assign SYNC = !I_1889_D;
  assign RED = I_67_S;
  assign GREEN = I_448_D;
  assign BLUE = I_768_D;
  assign I_1039_D = !(!I_3015_D && I_3499_D);
  assign I_1089_D = !(I_2371_S && !I_1731_D);
  assign I_1091_D = !(!I_2049_D && !I_453_D);

  always @(*)
    if (I_1571_D)
      I_1093_D <= 1'b0;
    else if (I_715_D)
      I_1093_D <= !I_1095_D;

  always @(*)
    if (I_1571_D)
      I_1095_D <= 1'b1;
    else if (!I_715_D)
      I_1095_D <= I_2073_D;

  assign I_1103_D = !(!I_2535_D && !I_3499_D);
  assign I_1111_D = I_1593_D? D4:!I_1271_D;
  assign I_1115_D = !(!I_1269_D && I_1275_D);

  always @(*)
    if (CLK)
      I_1119_D <= !I_959_D;

  assign I_1185_D = !(I_2371_S && I_2275_D);
  assign I_1211_D = !(!I_317_D && !I_797_D && !I_479_D);
  assign I_1213_D = !(!I_317_D && !I_479_D && !I_797_D);
  assign I_1251_D = !(I_1091_D && !I_311_D);

  always @(*)
    if (I_1571_D)
      I_1253_D <= 1'b0;
    else if (I_715_D)
      I_1253_D <= !I_1255_D;

  always @(*)
    if (I_1571_D)
      I_1255_D <= 1'b1;
    else if (!I_715_D)
      I_1255_D <= I_2233_D;

  always @(*)
    if (I_1119_D)
      I_1257_D <= !I_1419_D;

  always @(*)
    if (!I_1119_D)
      I_1259_D <= !I_1257_D;

  assign I_1265_D = I_1999_D? !I_2071_S:I_2071_S;

  always @(*)
    if (I_479_D)
      I_1267_D <= !I_3585_D;

  always @(*)
    if (!I_479_D)
      I_1269_D <= !I_1267_D;

  always @(*)
    if (I_479_D)
      I_1271_D <= !I_1431_D;

  assign I_1275_D = !(I_797_D && !I_479_D);
  assign I_1279_D = I_1213_D? !I_1119_D:I_1119_D;
  assign I_128_D = !(I_1089_D || I_225_D);

  always @(*)
    if (I_1571_D)
      I_133_D <= 1'b1;
    else if (I_395_D)
      I_133_D <= !I_135_D;

  assign I_1359_D = !(I_3499_D && !I_3175_D);

  always @(*)
    if (I_1571_D)
      I_135_D <= 1'b0;
    else if (!I_395_D)
      I_135_D <= I_2073_D;

  always @(*)
    if (I_1571_D)
      I_1413_D <= 1'b0;
    else if (I_715_D)
      I_1413_D <= !I_1415_D;

  always @(*)
    if (I_1571_D)
      I_1415_D <= 1'b1;
    else if (!I_715_D)
      I_1415_D <= I_2393_D;

  always @(*)
    if (I_1435_D)
      I_1417_D <= D7;

  always @(*)
    if (!I_1435_D)
      I_1419_D <= !I_1417_D;

  assign I_1423_D = !(!I_3499_D && !I_2695_D);
  assign I_1425_S = I_2071_S && I_1999_D;

  always @(*)
    if (CLK)
      I_1427_D <= !I_1429_D;

  always @(*)
    if (!CLK)
      I_1429_D <= !I_797_D;

  always @(*)
    if (!I_479_D)
      I_1431_D <= I_1433_D;

  assign I_1433_D = I_1593_D? D3:!I_953_D;
  assign I_1435_D = !(!I_317_D || I_797_D || !I_1119_D);

  always @(*)
    if (CLK)
      I_1439_D <= I_1439_S;

  assign I_1439_S = !(I_959_D && I_319_D && I_637_D);
  assign I_1499_D = !(!I_317_D && I_3499_D);
  assign I_1518_D = !(I_1359_D && I_1423_D);
  assign I_1535_D = !(I_1499_D && I_1119_D && I_3667_D);

  always @(*)
    if (!I_479_D)
      I_153_D <= I_155_D;

  assign I_155_D = I_1593_D? D0:1'b0;

  always @(*)
    if (I_1735_D)
      I_1569_D <= I_1891_S;

  always @(*)
    if (!I_1735_D)
      I_1571_D <= !I_1569_D;

  always @(*)
    if (!I_317_D)
      I_1573_D <= I_1575_D;

  always @(*)
    if (I_317_D)
      I_1575_D <= !I_1573_D;

  always @(*)
    if (!CLK)
      I_157_D <= I_1439_D && I_477_D;

  assign I_1585_D = !(I_1518_D && I_1679_D);

  always @(*)
    if (!CLK)
      I_1591_D <= I_1845_D;

  always @(*)
    if (CLK)
      I_1593_D <= !I_1591_D;

  assign I_1648_D = !(I_1518_D || I_1679_D);
  assign I_1673_D = !(!I_1251_D && !I_1259_D);
  assign I_1679_D = !(I_1743_D && I_1807_D);
  assign I_1693_D = !(I_1535_D && I_1695_D && I_1855_D);
  assign I_1695_D = !(I_1499_D && A11 && !I_1119_D);

  always @(*)
    if (I_1119_D)
      I_1729_D <= I_2275_D;

  always @(*)
    if (!I_1119_D)
      I_1731_D <= !I_1729_D;

  always @(*)
    if (!I_1575_D)
      I_1733_D <= I_1735_D;

  always @(*)
    if (I_1575_D)
      I_1735_D <= !I_1733_D;

  assign I_1737_D = !(!I_1259_D && I_1251_D);
  assign I_1743_D = !(!I_3015_D && !I_3499_D);
  assign I_1807_D = !(I_3499_D && !I_3495_D);
  assign I_1832_D = !(I_1673_D && I_1737_D);
  assign I_1845_D = !(!I_317_D && !I_797_D && I_457_D);
  assign I_1855_D = !(!I_1499_D && I_1119_D && I_1901_D);
  assign I_1889_D = !(!I_1571_D && I_1987_D);
  assign I_1891_S = !(I_1895_D && I_2055_D && !I_2215_D && !I_2375_D);

  always @(*)
    if (!I_1735_D)
      I_1893_D <= I_1895_D;

  always @(*)
    if (I_1735_D)
      I_1895_D <= !I_1893_D;

  assign I_1899_S = !(I_133_D || I_777_D);
  assign I_1901_D = !(I_133_D && !I_777_D);

  always @(*)
    if (!CLK)
      I_1911_D <= !I_1913_D;

  always @(*)
    if (CLK)
      I_1913_D <= I_1913_S;

  assign I_1913_S = !(!I_797_D || !I_479_D);
  assign I_1915_S = !(I_1119_D || I_1911_D);
  assign I_1917_D = !(I_1693_D && I_1911_D);
  assign I_1962_D = (!I_133_D || !I_777_D) && !I_1899_S;
  assign I_1987_D = !(I_2051_D && I_2115_D);
  assign I_1999_D = !(I_2063_D && I_2127_D);
  assign I_2011_D = !(I_2075_D && I_2139_D);
  assign I_2013_D = !(!I_1911_D && I_2011_D);
  assign I_2015_D = !(I_1499_D && I_1119_D && I_3669_D);

  always @(*)
    if (I_2369_D)
      I_2049_D <= !I_2209_D;

  assign I_2051_D = !(I_3075_D && !I_937_D);

  always @(*)
    if (!I_1895_D)
      I_2053_D <= I_2055_D;

  always @(*)
    if (I_1895_D)
      I_2055_D <= !I_2053_D;

  assign I_2063_D = !(!I_2855_D && !I_3499_D);
  assign I_2065_S = !(I_1585_D && !I_1648_D);
  assign I_2069_D = !(I_1518_D && !I_2215_D);
  assign I_2071_D = I_2055_D? I_2071_S:!I_2071_S;
  assign I_2071_S = !(I_1039_D && I_1103_D);

  always @(*)
    if (I_1435_D)
      I_2073_D <= D0;

  assign I_2075_D = !(I_2071_D && I_1499_D);
  assign I_2077_D = !(I_1917_D && I_2013_D);
  assign I_2115_D = !(I_937_D && !I_3491_S);
  assign I_2127_D = !(I_3499_D && !I_3335_D);
  assign I_2132_D = !(I_1518_D || !I_2215_D);
  assign I_2139_D = !(!I_1499_D && I_2073_D);
  assign I_2154_D = !(!I_2699_D || I_2539_S || I_3562_D);
  assign I_2173_D = !(I_2015_D && I_2175_D && I_2335_D);
  assign I_2175_D = !(I_1499_D && !I_1119_D && A12);

  always @(*)
    if (!I_2369_D)
      I_2209_D <= I_2049_D;

  assign I_2211_D = !(I_2055_D && I_2215_D);

  always @(*)
    if (!I_2055_D)
      I_2213_D <= I_2215_D;

  always @(*)
    if (I_2055_D)
      I_2215_D <= !I_2213_D;

  assign I_2225_D = !(I_1999_D && I_2319_D);
  assign I_2231_S = I_2071_S && !I_2055_D;

  always @(*)
    if (I_1435_D)
      I_2233_D <= D1;

  assign I_2235_D = !(I_1499_D && I_2549_D);
  assign I_2237_D = !(I_2173_D && I_1911_D);
  assign I_225_D = !I_1832_D && !I_227_D || !I_289_D;
  assign I_2275_D = !(I_2211_D && !I_2375_D);
  assign I_227_D = !(I_291_D && I_355_D);
  assign I_2288_D = !(I_1999_D || I_2319_D);
  assign I_2319_D = !(I_2383_D && I_2447_D);
  assign I_2331_D = !(!I_1499_D && I_2233_D);
  assign I_2333_D = !(!I_1911_D && I_2395_D);
  assign I_2335_D = !(!I_1499_D && I_1119_D);
  assign I_235_D = !(I_2553_D && I_2713_D && !I_553_D);

  always @(*)
    if (I_2689_D)
      I_2369_D <= !I_2529_D;

  assign I_2371_S = !(!I_3815_D || I_2632_D);

  always @(*)
    if (!I_2215_D)
      I_2373_D <= I_2375_D;

  always @(*)
    if (I_2215_D)
      I_2375_D <= !I_2373_D;

  assign I_2379_S = !(I_3337_D || I_3499_D);
  assign I_2383_D = !(!I_3499_D && !I_3175_D);
  assign I_2391_D = !(I_1265_D && !I_2375_D);

  always @(*)
    if (I_1435_D)
      I_2393_D <= D2;

  assign I_2395_D = !(I_2235_D && I_2331_D);
  assign I_2397_D = !(I_2237_D && I_2333_D);
  assign I_2447_D = !(I_3499_D && I_3337_D);
  assign I_2454_D = !(I_1265_D || !I_2375_D);
  assign I_2491_D = !(!I_1499_D && I_2393_D);
  assign I_2493_D = !(!I_1911_D && I_2650_D);
  assign I_2495_D = !(I_1499_D && I_1119_D && !I_3829_S);

  always @(*)
    if (!I_2689_D)
      I_2529_D <= I_2369_D;

  always @(*)
    if (I_3177_D)
      I_2533_D <= 1'b0;
    else if (!I_1571_D)
      I_2533_D <= I_2535_D;

  always @(*)
    if (I_3177_D)
      I_2535_D <= 1'b1;
    else if (I_1571_D)
      I_2535_D <= !I_2533_D;

  assign I_2539_S = !(!I_3655_D || !I_3815_D);
  assign I_2545_S = !I_1585_D || !I_1648_D && I_1425_S;
  assign I_2549_D = I_2231_S? I_2549_S:!I_2549_S;
  assign I_2549_S = !(I_2069_D && !I_2132_D);

  always @(*)
    if (I_1435_D)
      I_2553_D <= D3;

  assign I_2555_D = !(I_1499_D && I_2871_D);
  assign I_2557_D = !(I_1911_D && I_2653_D);
  assign I_2632_D = !(I_3335_D || I_3495_D || I_3655_D);
  assign I_2634_D = !(I_3495_D || I_3655_D || !I_3815_D);
  assign I_2650_D = !(I_2491_D && I_2555_D);
  assign I_2653_D = !(I_2495_D && I_2655_D && I_2815_D);
  assign I_2655_D = !(I_1499_D && !I_1119_D && A13);

  always @(*)
    if (I_3009_D)
      I_2689_D <= !I_2849_D;

  always @(*)
    if (I_3177_D)
      I_2693_D <= 1'b0;
    else if (!I_2535_D)
      I_2693_D <= I_2695_D;

  always @(*)
    if (I_3177_D)
      I_2695_D <= 1'b1;
    else if (I_2535_D)
      I_2695_D <= !I_2693_D;

  assign I_2699_D = !(I_2634_D && I_2794_D);
  assign I_2705_S = !(I_2225_D && !I_2288_D);
  assign I_2709_D = I_2869_D? !I_2709_S:I_2709_S;
  assign I_2709_S = I_1425_S? I_2065_S:!I_2065_S;
  assign I_2711_S = !I_2069_D || !I_2132_D && I_2231_S;

  always @(*)
    if (I_1435_D)
      I_2713_D <= D4;

  assign I_2715_D = !(I_2709_D && I_1499_D);
  assign I_2717_D = !(I_2493_D && I_2557_D);
  assign I_2794_D = !(!I_3015_D || !I_3175_D || !I_3335_D);
  assign I_2811_D = !(!I_1499_D && I_2553_D);
  assign I_2813_D = !(!I_1911_D && I_2875_D);
  assign I_2815_D = !(!I_777_D && !I_1499_D && I_1119_D);

  always @(*)
    if (!I_3009_D)
      I_2849_D <= I_2689_D;

  always @(*)
    if (I_3177_D)
      I_2853_D <= 1'b0;
    else if (!I_2695_D)
      I_2853_D <= I_2855_D;

  always @(*)
    if (I_3177_D)
      I_2855_D <= 1'b1;
    else if (I_2695_D)
      I_2855_D <= !I_2853_D;

  assign I_2865_D = !(I_1679_D && I_3116_D);
  assign I_2869_D = !I_2391_D || !I_2454_D && I_2711_S;
  assign I_2871_D = I_2711_S? I_2871_S:!I_2871_S;
  assign I_2871_S = !(I_2391_D && !I_2454_D);

  always @(*)
    if (I_1435_D)
      I_2873_D <= D5;

  assign I_2875_D = !(I_2715_D && I_2811_D);
  assign I_2877_D = !(I_1911_D && I_3133_D);
  assign I_289_D = !(I_1832_D && I_227_D);
  assign I_291_D = !(I_1251_D && !I_613_D);
  assign I_2928_D = !(I_1679_D || I_3116_D);

  always @(*)
    if (I_1571_D)
      I_293_D <= 1'b1;
    else if (I_395_D)
      I_293_D <= !I_295_D;

  assign I_2953_D = !(I_937_D && I_2955_D);
  assign I_2955_D = !(!I_3015_D && !I_3175_D && !I_3335_D && !I_3815_D);
  assign I_2957_D = !(I_3499_D && I_3339_D);

  always @(*)
    if (I_1571_D)
      I_295_D <= 1'b0;
    else if (!I_395_D)
      I_295_D <= I_2233_D;

  assign I_2971_D = !(!I_1499_D && I_2713_D);
  assign I_2972_D = !(I_2813_D && I_2877_D);
  assign I_2975_D = !(I_3829_S && I_1499_D && I_1119_D);

  always @(*)
    if (I_3329_D)
      I_3009_D <= !I_3169_D;

  always @(*)
    if (I_3177_D)
      I_3013_D <= 1'b0;
    else if (!I_2855_D)
      I_3013_D <= I_3015_D;

  always @(*)
    if (I_3177_D)
      I_3015_D <= 1'b1;
    else if (I_2855_D)
      I_3015_D <= !I_3013_D;

  assign I_3017_D = !(!I_937_D && I_3083_D);
  assign I_3021_D = !(!I_3499_D && !I_3335_D);
  assign I_3023_D = !(!I_2379_S && I_3116_D);
  assign I_3027_D = I_3189_S? !I_3985_D:I_3985_D;
  assign I_3029_D = I_3191_S? !I_3345_D:I_3345_D;
  assign I_3031_D = I_3191_D? !I_3031_S:I_3031_S;
  assign I_3031_S = I_2545_S? I_2705_S:!I_2705_S;

  always @(*)
    if (I_1435_D)
      I_3033_D <= D6;

  assign I_3035_D = !(I_1499_D && I_3031_D);
  assign I_3075_D = !(I_2632_D && !I_2855_D && I_3171_D && I_3175_D);
  assign I_3083_D = !(!I_3015_D && !I_3815_D);
  assign I_3086_D = !(!I_2379_S || I_3116_D);
  assign I_3112_D = !(I_2953_D && I_3017_D);
  assign I_3116_D = !(I_2957_D && I_3021_D);

  always @(*)
    if (I_479_D)
      I_311_D <= !I_471_D;

  assign I_3130_D = !(I_2971_D && I_3035_D);
  assign I_3133_D = !(I_2975_D && I_3135_D);
  assign I_3135_D = !(I_1499_D && !I_1119_D && A14);

  always @(*)
    if (I_479_D)
      I_313_D <= !I_153_D;

  always @(*)
    if (!I_3329_D)
      I_3169_D <= I_3009_D;

  assign I_3171_D = !(I_3015_D && I_3175_D);

  always @(*)
    if (I_3177_D)
      I_3173_D <= 1'b0;
    else if (!I_3015_D)
      I_3173_D <= I_3175_D;

  always @(*)
    if (I_3177_D)
      I_3175_D <= 1'b1;
    else if (I_3015_D)
      I_3175_D <= !I_3173_D;

  assign I_3177_D = !I_3112_D;

  always @(*)
    if (CLK)
      I_317_D <= !I_157_D;

  assign I_3185_S = !I_2225_D || !I_2288_D && I_2545_S;
  assign I_3189_S = I_3345_D && I_3191_S;
  assign I_3191_D = I_2709_S && I_2869_D;
  assign I_3191_S = I_3031_S && I_3191_D;
  assign I_3193_D = !(I_1911_D && I_3449_D);
  assign I_3197_D = !(I_1911_D && I_3453_D);

  always @(*)
    if (!CLK)
      I_319_D <= I_1439_D && I_479_D;

  assign I_3285_D = !(I_3349_D && I_3413_D);
  assign I_3287_D = !(I_3347_D && I_1499_D && I_1119_D);
  assign I_3289_D = !(!I_1911_D && I_3285_D);
  assign I_3291_D = !(I_1499_D && I_1119_D);
  assign I_3293_D = !(!I_1911_D && I_3130_D);

  always @(*)
    if (I_3815_D)
      I_3329_D <= !I_3489_D;

  always @(*)
    if (!I_3112_D)
      I_3333_D <= 1'b0;
    else if (!I_3175_D)
      I_3333_D <= I_3335_D;

  always @(*)
    if (!I_3112_D)
      I_3335_D <= 1'b1;
    else if (I_3175_D)
      I_3335_D <= !I_3333_D;

  assign I_3337_D = I_3655_D? I_3499_D:!I_3499_D;
  assign I_3339_D = I_3499_D? !I_3497_S:I_3497_S;
  assign I_3345_D = I_3185_S? I_3345_S:!I_3345_S;
  assign I_3345_S = !(I_2865_D && !I_2928_D);
  assign I_3347_D = I_3507_D? !I_3503_D:I_3503_D;
  assign I_3349_D = !(!I_1895_D && I_1499_D);
  assign I_3353_D = !(I_3193_D && I_3289_D);
  assign I_3357_D = !(I_3197_D && I_3293_D);
  assign I_3413_D = !(I_3906_D && !I_1499_D);
  assign I_3427_D = !(I_2855_D && I_3015_D);
  assign I_3447_D = !(I_1499_D && !I_1119_D && A10);
  assign I_3449_D = !(I_3287_D && I_3447_D && I_3607_D);
  assign I_3451_D = !(I_1499_D && !I_1119_D && A15);
  assign I_3453_D = !(I_3291_D && I_3451_D && I_3611_D);

  always @(*)
    if (!I_3815_D)
      I_3489_D <= I_3329_D;

  assign I_3491_S = !(I_3427_D || I_3587_D);

  always @(*)
    if (!I_3112_D)
      I_3493_D <= 1'b0;
    else if (!I_3335_D)
      I_3493_D <= I_3495_D;

  always @(*)
    if (!I_3112_D)
      I_3495_D <= 1'b1;
    else if (I_3335_D)
      I_3495_D <= !I_3493_D;

  assign I_3497_S = I_3499_D && !I_3655_D;
  assign I_3499_D = !(!I_2154_D && I_777_D);
  assign I_3499_S = I_3497_S && I_3499_D;
  assign I_3501_D = !(!I_3495_D && !I_3499_D);
  assign I_3503_D = I_3825_D? I_3503_S:!I_3503_S;
  assign I_3503_S = !(I_3023_D && !I_3086_D);
  assign I_3505_D = !(I_2319_D && I_3663_S);
  assign I_3507_D = I_3985_D && I_3189_S;
  assign I_3517_D = !(I_1911_D && I_3773_D);
  assign I_355_D = !(!I_1093_D && !I_1251_D);
  assign I_3562_D = !(!I_3495_D || !I_3815_D);
  assign I_3565_D = !(I_3499_D && I_3499_S);
  assign I_3568_D = !(I_2319_D || I_3663_S);
  assign I_3585_D = !(I_3913_S && I_3975_D);
  assign I_3587_D = !(I_3175_D && I_3335_D && !I_3815_D);
  assign I_3607_D = !(I_1962_D && !I_1499_D && I_1119_D);
  assign I_3609_D = !(I_3027_D && I_1499_D && I_1119_D);
  assign I_3611_D = !(!I_1499_D && I_1119_D);
  assign I_3613_D = !(!I_1911_D && I_3997_D);
  assign I_3615_D = !(I_3029_D && I_1499_D && I_1119_D);

  always @(*)
    if (!I_3112_D)
      I_3653_D <= 1'b0;
    else if (!I_3495_D)
      I_3653_D <= I_3655_D;

  always @(*)
    if (!I_3112_D)
      I_3655_D <= 1'b1;
    else if (I_3495_D)
      I_3655_D <= !I_3653_D;

  assign I_3663_D = I_3823_D? !I_3663_S:I_3663_S;
  assign I_3663_S = !(I_3501_D && I_3565_D);
  assign I_3667_D = I_3827_D? !I_3663_D:I_3663_D;
  assign I_3669_D = I_3829_D? !I_3669_S:I_3669_S;
  assign I_3669_S = I_3823_S? I_2379_S:!I_2379_S;
  assign I_3677_D = !(I_3517_D && I_3613_D);
  assign I_3725_D = !(!A13 && !A14 && !A12 && !A15);
  assign I_3745_D = !(!I_2855_D && !I_293_D);
  assign I_3747_D = !(!I_3015_D && !I_293_D);
  assign I_3753_D = !(I_3453_D && I_3133_D && !nMAP);
  assign I_3755_S = !(I_3725_D || I_3883_D);
  assign I_3767_D = !(!I_1499_D && I_3904_D);
  assign I_3769_D = !(I_1499_D && !I_1119_D && A9);
  assign I_3771_D = !(I_3609_D && I_3769_D && I_3929_D);
  assign I_3773_D = !(I_3615_D && I_3775_D && I_3935_D);
  assign I_3775_D = !(I_1499_D && !I_1119_D && A8);
  assign I_3809_D = !(!I_2695_D && I_293_D);
  assign I_3811_D = !(!I_2855_D && I_293_D);

  always @(*)
    if (!I_3112_D)
      I_3813_D <= 1'b0;
    else if (!I_3655_D)
      I_3813_D <= I_3815_D;

  always @(*)
    if (!I_3112_D)
      I_3815_D <= 1'b1;
    else if (I_3655_D)
      I_3815_D <= !I_3813_D;

  assign I_3817_D = !(!I_3453_D && nMAP);
  assign I_3823_D = !I_3023_D || !I_3086_D && I_3825_D;
  assign I_3823_S = I_3663_S && I_3823_D;
  assign I_3825_D = !I_3505_D || !I_3568_D && I_3825_S;
  assign I_3825_S = !I_2865_D || !I_2928_D && I_3185_S;
  assign I_3827_D = I_3503_D && I_3507_D;
  assign I_3829_D = I_3663_D && I_3827_D;
  assign I_3829_S = I_3669_S && I_3829_D;
  assign I_3831_D = !(I_1499_D && !I_1735_D);
  assign I_3835_D = !(I_3771_D && I_1911_D);
  assign I_3837_D = !(!I_1575_D && I_1499_D);
  assign I_3883_D = !(!A11 && A9 && !A10 && A8);
  assign I_3884_D = !(RnW && A14 && nMAP && A15);
  assign I_3904_D = !(I_3745_D && I_3809_D);
  assign I_3906_D = !(I_3747_D && I_3811_D);
  assign I_3909_D = !(!I_2695_D && !I_293_D);
  assign I_3911_D = !(I_293_D && !I_2535_D);
  assign I_3913_S = !(I_3753_D && I_3817_D && I_3977_D);
  assign I_3926_D = !(I_3767_D && I_3831_D);
  assign I_3929_D = !(I_3033_D && !I_1499_D && I_1119_D);
  assign I_3931_D = !(!I_1911_D && I_3926_D);
  assign I_3933_D = !(!I_1499_D && I_3973_D);
  assign I_3935_D = !(I_2873_D && !I_1499_D && I_1119_D);
  assign I_395_D = !(I_2553_D && !I_2713_D && !I_553_D);
  assign I_3973_D = !(I_3909_D && I_3911_D);
  assign I_3975_D = !(I_3755_S && !I_1119_D);
  assign I_3977_D = !(!I_3133_D && nMAP);
  assign I_3981_D = !(!RnW && !I_1119_D);
  assign I_3985_D = I_3825_S? I_3985_S:!I_3985_S;
  assign I_3985_S = !(I_3505_D && !I_3568_D);
  assign I_3995_D = !(I_3835_D && I_3931_D);
  assign I_3997_D = !(I_3837_D && I_3933_D);
  assign I_448_D = !(I_1089_D || I_545_D);

  always @(*)
    if (I_1571_D)
      I_453_D <= 1'b1;
    else if (I_395_D)
      I_453_D <= !I_455_D;

  always @(*)
    if (I_1571_D)
      I_455_D <= 1'b0;
    else if (!I_395_D)
      I_455_D <= I_2393_D;

  assign I_457_D = !(!I_2873_D && !I_3033_D);

  always @(*)
    if (!I_479_D)
      I_471_D <= I_631_D;

  always @(*)
    if (!I_479_D)
      I_473_D <= I_475_D;

  assign I_475_D = I_1593_D? D1:!I_313_D;
  assign I_477_D = I_573_D? !I_317_D:I_317_D;

  always @(*)
    if (CLK)
      I_479_D <= !I_319_D;

  assign I_524_D = !(I_1211_D || I_1185_D);
  assign I_545_D = !I_1832_D && !I_547_D || !I_609_D;
  assign I_547_D = !(I_611_D && I_675_D);
  assign I_553_D = !(!I_2873_D && !I_3033_D && I_524_D);
  assign I_555_D = !(I_2713_D && !I_2553_D && !I_553_D);
  assign I_573_D = !(!I_479_D && !I_797_D);
  assign I_609_D = !(I_1832_D && I_547_D);
  assign I_611_D = !(I_1251_D && !I_773_D);

  always @(*)
    if (I_1571_D)
      I_613_D <= 1'b1;
    else if (I_555_D)
      I_613_D <= !I_615_D;

  always @(*)
    if (I_1571_D)
      I_615_D <= 1'b0;
    else if (!I_555_D)
      I_615_D <= I_2073_D;

  assign I_631_D = I_1593_D? D5:!I_791_D;

  always @(*)
    if (I_479_D)
      I_633_D <= !I_473_D;

  always @(*)
    if (!CLK)
      I_637_D <= I_1439_D && I_957_D;

  assign I_675_D = !(!I_1253_D && !I_1251_D);
  assign I_67_S = !(I_1889_D || !I_128_D);
  assign I_715_D = !(!I_2713_D && !I_2553_D && !I_553_D);
  assign I_768_D = !(I_1089_D || I_865_D);

  always @(*)
    if (I_1571_D)
      I_773_D <= 1'b1;
    else if (I_555_D)
      I_773_D <= !I_775_D;

  always @(*)
    if (I_1571_D)
      I_775_D <= 1'b0;
    else if (!I_555_D)
      I_775_D <= I_2233_D;

  always @(*)
    if (!I_235_D)
      I_777_D <= I_2393_D;

  always @(*)
    if (I_479_D)
      I_791_D <= !I_951_D;

  always @(*)
    if (!I_479_D)
      I_793_D <= I_795_D;

  assign I_795_D = I_1593_D? D2:!I_633_D;

  always @(*)
    if (CLK)
      I_797_D <= !I_637_D;

  assign I_865_D = !I_1832_D && !I_867_D || !I_929_D;
  assign I_867_D = !(I_931_D && I_995_D);
  assign I_929_D = !(I_1832_D && I_867_D);
  assign I_931_D = !(I_1251_D && !I_933_D);

  always @(*)
    if (I_1571_D)
      I_933_D <= 1'b1;
    else if (I_555_D)
      I_933_D <= !I_935_D;

  always @(*)
    if (I_1571_D)
      I_935_D <= 1'b0;
    else if (!I_555_D)
      I_935_D <= I_2393_D;

  always @(*)
    if (!I_235_D)
      I_937_D <= I_2233_D;

  always @(*)
    if (!I_479_D)
      I_951_D <= I_1111_D;

  always @(*)
    if (I_479_D)
      I_953_D <= !I_793_D;

  assign I_957_D = I_479_D? !I_797_D:I_797_D;

  always @(*)
    if (!CLK)
      I_959_D <= I_1439_D && I_1279_D;

  assign I_995_D = !(!I_1251_D && !I_1413_D);

endmodule
