//----------------------------------------------------------------------------
//
//  ORIC ULA Verilog CMOS netlist
//
//  Erik Persson, 2023
//
//  Building on earlier work by Lance Ewing, Mike Connors and Mike Brown
//
//  Changelog
//  - Started with file 001_top_unprocessed.v
//  - Added ports, guided by 006_mjb_sorted.v
//  - Dos2unix and tab => 2 spaces
//  - Repaired nets based on comments in 006_mjb_sorted.v
//
//----------------------------------------------------------------------------

module Top
(
  input  supply1 VDD,   // Positive voltage
  input  supply0 VSS,   // Ground

  input  wire    CLK,   // 12 MHz clock

  // 6502 Address bus high byte
  input  wire    A8,
  input  wire    A9,
  input  wire    A10,
  input  wire    A11,
  input  wire    A12,
  input  wire    A13,
  input  wire    A14,
  input  wire    A15,

  // 6502 data bus
  input  wire    D0,
  input  wire    D1,
  input  wire    D2,
  input  wire    D3,
  input  wire    D4,
  input  wire    D5,
  input  wire    D6,
  input  wire    D7,

  input  wire    RnW,    // 6502 read cycle indicator
  input  wire    nMAP,   // From expansion bus

  // DRAM Row and column address
  output wire    RC0,
  output wire    RC1,
  output wire    RC2,
  output wire    RC3,
  output wire    RC4,
  output wire    RC5,
  output wire    RC6,
  output wire    RC7,

  output wire    MXSEL,   // DRAM mux select
  output wire    nROM,    // ROM chip select
  output wire    PHI,     // Output clock
  output wire    CAS,     // DRAM Column Access Strobe, active high
  output wire    RAS,     // DRAM Row Access Strobe, active high
  output wire    WE,      // DRAM Write Enable, active high
  output wire    nIO,     // 6522 chip select

  output wire    SYNC,    // Composite sync signal
  output wire    RED,     // Red video output
  output wire    GREEN,   // Green video output
  output wire    BLUE     // Blue video output
);

wire  I_1002_D;
wire  I_1003_D;
wire  I_1003_G;
wire  I_1004_D;
wire  I_1005_D;
wire  I_1005_G;
wire  I_1008_D;
wire  I_1009_D;
wire  I_1009_G;
wire  I_1010_D;
wire  I_1011_D;
wire  I_1011_G;
wire  I_1014_D;
wire  I_1015_D;
wire  I_1019_G;
wire  I_101_D;
wire  I_1022_D;
wire  I_1025_D;
wire  I_1025_G;
wire  I_1027_S;
wire  I_1028_D;
wire  I_1029_D;
wire  I_1033_D;
wire  I_1034_D;
wire  I_1034_S;
wire  I_1035_D;
wire  I_1035_G;
wire  I_1035_S;
wire  I_1036_D;
wire  I_1036_S;
wire  I_1037_D;
wire  I_1037_G;
wire  I_1037_S;
wire  I_1038_D;
wire  I_1039_D;
wire  I_103_D;
wire  I_1040_D;
wire  I_1040_S;
wire  I_1041_D;
wire  I_1041_G;
wire  I_1041_S;
wire  I_1042_D;
wire  I_1042_S;
wire  I_1043_D;
wire  I_1043_G;
wire  I_1043_S;
wire  I_1045_D;
wire  I_1046_S;
wire  I_1047_G;
wire  I_1047_S;
wire  I_1049_S;
wire  I_104_D;
wire  I_104_G;
wire  I_1051_S;
wire  I_1055_S;
wire  I_105_D;
wire  I_1061_D;
wire  I_1063_D;
wire  I_1065_D;
wire  I_1067_D;
wire  I_1069_D;
wire  I_106_D;
wire  I_106_G;
wire  I_1072_D;
wire  I_1072_G;
wire  I_1073_D;
wire  I_1074_D;
wire  I_1074_G;
wire  I_1075_D;
wire  I_1076_D;
wire  I_1076_G;
wire  I_1077_D;
wire  I_107_D;
wire  I_1085_D;
wire  I_1087_D;
wire  I_1088_D;
wire  I_1089_D;
wire  I_108_D;
wire  I_108_G;
wire  I_1090_D;
wire  I_1091_D;
wire  I_1093_D;
wire  I_1093_S;
wire  I_1095_D;
wire  I_1096_G;
wire  I_1096_S;
wire  I_1097_S;
wire  I_1098_G;
wire  I_1098_S;
wire  I_1099_S;
wire  I_109_D;
wire  I_10_D;
wire  I_1100_G;
wire  I_1100_S;
wire  I_1101_S;
wire  I_1102_D;
wire  I_1103_D;
wire  I_1104_D;
wire  I_1104_G;
wire  I_1104_S;
wire  I_1105_D;
wire  I_1105_G;
wire  I_1105_S;
wire  I_1106_D;
wire  I_1106_G;
wire  I_1106_S;
wire  I_1107_D;
wire  I_1107_G;
wire  I_1107_S;
wire  I_1108_D;
wire  I_1108_G;
wire  I_1108_S;
wire  I_1109_D;
wire  I_1109_G;
wire  I_1109_S;
wire  I_110_D;
wire  I_110_G;
wire  I_1111_D;
wire  I_1112_D;
wire  I_1113_D;
wire  I_1113_S;
wire  I_1114_D;
wire  I_1115_D;
wire  I_1116_G;
wire  I_1116_S;
wire  I_1117_D;
wire  I_1119_D;
wire  I_111_D;
wire  I_1120_D;
wire  I_1121_D;
wire  I_1121_G;
wire  I_112_D;
wire  I_112_G;
wire  I_1132_D;
wire  I_1133_D;
wire  I_1133_G;
wire  I_1136_D;
wire  I_1137_D;
wire  I_1137_G;
wire  I_1139_D;
wire  I_113_D;
wire  I_1144_D;
wire  I_1145_D;
wire  I_1145_G;
wire  I_114_D;
wire  I_114_G;
wire  I_1153_G;
wire  I_1158_D;
wire  I_115_D;
wire  I_1164_D;
wire  I_1165_D;
wire  I_1165_G;
wire  I_1166_D;
wire  I_1168_D;
wire  I_1169_D;
wire  I_1169_G;
wire  I_116_D;
wire  I_116_G;
wire  I_1178_D;
wire  I_117_D;
wire  I_1180_D;
wire  I_1183_G;
wire  I_1184_D;
wire  I_1185_D;
wire  I_1185_G;
wire  I_1187_S;
wire  I_1188_D;
wire  I_1189_D;
wire  I_118_D;
wire  I_118_G;
wire  I_1193_G;
wire  I_1195_D;
wire  I_1196_D;
wire  I_1196_S;
wire  I_1197_D;
wire  I_1197_G;
wire  I_1197_S;
wire  I_1198_S;
wire  I_1199_G;
wire  I_1199_S;
wire  I_11_D;
wire  I_11_G;
wire  I_1200_D;
wire  I_1200_S;
wire  I_1201_D;
wire  I_1201_G;
wire  I_1201_S;
wire  I_1205_D;
wire  I_1207_D;
wire  I_1208_D;
wire  I_1209_D;
wire  I_1209_S;
wire  I_1210_D;
wire  I_1211_D;
wire  I_1212_D;
wire  I_1213_D;
wire  I_1221_D;
wire  I_1223_D;
wire  I_1225_D;
wire  I_1227_D;
wire  I_1228_D;
wire  I_1228_G;
wire  I_1230_D;
wire  I_1230_G;
wire  I_1235_D;
wire  I_1237_D;
wire  I_1239_D;
wire  I_1244_D;
wire  I_1244_G;
wire  I_1247_D;
wire  I_1249_D;
wire  I_1250_D;
wire  I_1250_G;
wire  I_1251_D;
wire  I_1253_D;
wire  I_1253_S;
wire  I_1255_D;
wire  I_1257_D;
wire  I_1258_G;
wire  I_1259_D;
wire  I_1259_S;
wire  I_1260_G;
wire  I_1261_G;
wire  I_1261_S;
wire  I_1262_G;
wire  I_1263_G;
wire  I_1263_S;
wire  I_1265_D;
wire  I_1267_D;
wire  I_1267_S;
wire  I_1269_D;
wire  I_1269_S;
wire  I_1271_D;
wire  I_1272_D;
wire  I_1273_D;
wire  I_1273_S;
wire  I_1274_D;
wire  I_1275_D;
wire  I_1279_D;
wire  I_1279_S;
wire  I_127_D;
wire  I_1280_D;
wire  I_1281_D;
wire  I_1281_G;
wire  I_1283_D;
wire  I_128_D;
wire  I_1292_D;
wire  I_1293_D;
wire  I_1293_G;
wire  I_1295_D;
wire  I_1297_D;
wire  I_1298_D;
wire  I_1299_D;
wire  I_1299_G;
wire  I_129_D;
wire  I_12_D;
wire  I_1301_D;
wire  I_1304_D;
wire  I_1305_D;
wire  I_1305_G;
wire  I_1307_D;
wire  I_1309_D;
wire  I_130_G;
wire  I_130_S;
wire  I_1311_G;
wire  I_1313_G;
wire  I_1318_D;
wire  I_131_S;
wire  I_1324_D;
wire  I_1325_D;
wire  I_1325_G;
wire  I_1329_G;
wire  I_1331_D;
wire  I_1335_D;
wire  I_133_D;
wire  I_133_S;
wire  I_1340_D;
wire  I_1341_D;
wire  I_1342_D;
wire  I_1343_D;
wire  I_1344_D;
wire  I_1345_D;
wire  I_1347_D;
wire  I_1348_D;
wire  I_1349_D;
wire  I_1355_D;
wire  I_1356_D;
wire  I_1356_S;
wire  I_1357_D;
wire  I_1357_G;
wire  I_1357_S;
wire  I_1358_D;
wire  I_1359_D;
wire  I_135_D;
wire  I_1361_S;
wire  I_1362_D;
wire  I_1363_D;
wire  I_1364_D;
wire  I_1365_D;
wire  I_1365_S;
wire  I_1368_D;
wire  I_1369_D;
wire  I_1369_S;
wire  I_136_D;
wire  I_136_G;
wire  I_136_S;
wire  I_1371_D;
wire  I_1373_S;
wire  I_1374_S;
wire  I_1375_G;
wire  I_1375_S;
wire  I_1379_D;
wire  I_137_D;
wire  I_137_G;
wire  I_137_S;
wire  I_1381_D;
wire  I_1383_D;
wire  I_1385_D;
wire  I_1387_D;
wire  I_1388_D;
wire  I_1388_G;
wire  I_138_D;
wire  I_138_G;
wire  I_138_S;
wire  I_1393_D;
wire  I_1397_D;
wire  I_1399_D;
wire  I_139_D;
wire  I_139_G;
wire  I_139_S;
wire  I_13_D;
wire  I_13_G;
wire  I_1401_D;
wire  I_1402_D;
wire  I_1402_G;
wire  I_1403_D;
wire  I_1407_D;
wire  I_1408_D;
wire  I_1408_G;
wire  I_1409_D;
wire  I_1409_G;
wire  I_140_D;
wire  I_140_G;
wire  I_140_S;
wire  I_1410_G;
wire  I_1410_S;
wire  I_1411_S;
wire  I_1413_D;
wire  I_1413_S;
wire  I_1415_D;
wire  I_1415_S;
wire  I_1417_D;
wire  I_1417_S;
wire  I_1419_D;
wire  I_1419_S;
wire  I_141_D;
wire  I_141_G;
wire  I_141_S;
wire  I_1420_S;
wire  I_1421_G;
wire  I_1421_S;
wire  I_1422_D;
wire  I_1423_D;
wire  I_1425_S;
wire  I_1427_D;
wire  I_1429_D;
wire  I_142_D;
wire  I_142_G;
wire  I_142_S;
wire  I_1431_D;
wire  I_1433_D;
wire  I_1435_D;
wire  I_1435_G;
wire  I_1435_S;
wire  I_1437_D;
wire  I_1439_D;
wire  I_1439_S;
wire  I_143_D;
wire  I_143_G;
wire  I_143_S;
wire  I_1448_D;
wire  I_1449_D;
wire  I_1449_G;
wire  I_144_D;
wire  I_144_G;
wire  I_144_S;
wire  I_1452_D;
wire  I_1453_D;
wire  I_1453_G;
wire  I_1456_D;
wire  I_1457_D;
wire  I_1457_G;
wire  I_145_D;
wire  I_145_G;
wire  I_145_S;
wire  I_1461_D;
wire  I_1469_D;
wire  I_146_D;
wire  I_146_G;
wire  I_146_S;
wire  I_1478_D;
wire  I_147_D;
wire  I_147_G;
wire  I_147_S;
wire  I_1480_D;
wire  I_1481_D;
wire  I_1481_G;
wire  I_1482_D;
wire  I_1483_D;
wire  I_1484_D;
wire  I_1485_D;
wire  I_1485_G;
wire  I_1486_D;
wire  I_1488_D;
wire  I_1489_D;
wire  I_1489_G;
wire  I_148_D;
wire  I_148_G;
wire  I_148_S;
wire  I_1491_D;
wire  I_1498_D;
wire  I_1499_D;
wire  I_149_D;
wire  I_149_G;
wire  I_149_S;
wire  I_14_D;
wire  I_1502_D;
wire  I_1507_D;
wire  I_1508_D;
wire  I_1511_S;
wire  I_1512_D;
wire  I_1512_S;
wire  I_1513_D;
wire  I_1513_G;
wire  I_1513_S;
wire  I_1515_S;
wire  I_1516_D;
wire  I_1516_S;
wire  I_1517_D;
wire  I_1517_G;
wire  I_1517_S;
wire  I_1518_D;
wire  I_1518_S;
wire  I_1519_G;
wire  I_1519_S;
wire  I_151_D;
wire  I_151_G;
wire  I_1520_D;
wire  I_1520_S;
wire  I_1521_D;
wire  I_1521_G;
wire  I_1521_S;
wire  I_1523_S;
wire  I_1525_D;
wire  I_1529_D;
wire  I_1531_S;
wire  I_1534_D;
wire  I_1535_D;
wire  I_1537_D;
wire  I_1539_D;
wire  I_153_D;
wire  I_1541_D;
wire  I_1544_D;
wire  I_1544_G;
wire  I_1546_D;
wire  I_1546_G;
wire  I_1547_D;
wire  I_1548_D;
wire  I_1548_G;
wire  I_1549_D;
wire  I_1550_D;
wire  I_1550_G;
wire  I_1551_D;
wire  I_1554_D;
wire  I_1554_G;
wire  I_1555_D;
wire  I_1559_D;
wire  I_155_D;
wire  I_1561_D;
wire  I_1569_D;
wire  I_1571_D;
wire  I_1571_S;
wire  I_1573_D;
wire  I_1573_S;
wire  I_1575_D;
wire  I_1575_S;
wire  I_1576_S;
wire  I_1577_G;
wire  I_1577_S;
wire  I_1578_D;
wire  I_1578_G;
wire  I_1578_S;
wire  I_1579_D;
wire  I_1579_G;
wire  I_1579_S;
wire  I_157_D;
wire  I_1580_D;
wire  I_1580_G;
wire  I_1580_S;
wire  I_1581_D;
wire  I_1581_G;
wire  I_1581_S;
wire  I_1582_D;
wire  I_1582_G;
wire  I_1582_S;
wire  I_1583_D;
wire  I_1583_G;
wire  I_1583_S;
wire  I_1584_D;
wire  I_1585_D;
wire  I_1586_D;
wire  I_1586_G;
wire  I_1586_S;
wire  I_1587_D;
wire  I_1587_G;
wire  I_1587_S;
wire  I_1588_S;
wire  I_1589_S;
wire  I_158_G;
wire  I_158_S;
wire  I_1591_D;
wire  I_1593_D;
wire  I_1593_S;
wire  I_1597_D;
wire  I_1598_S;
wire  I_1599_S;
wire  I_159_S;
wire  I_15_D;
wire  I_15_G;
wire  I_1609_D;
wire  I_1610_D;
wire  I_1611_D;
wire  I_1611_G;
wire  I_1612_D;
wire  I_1613_D;
wire  I_1613_G;
wire  I_1614_D;
wire  I_1615_D;
wire  I_1615_G;
wire  I_1618_D;
wire  I_1619_D;
wire  I_1619_G;
wire  I_1620_D;
wire  I_1621_D;
wire  I_1621_G;
wire  I_1623_D;
wire  I_1627_D;
wire  I_162_D;
wire  I_1631_G;
wire  I_1638_D;
wire  I_163_D;
wire  I_163_G;
wire  I_1642_D;
wire  I_1643_D;
wire  I_1643_G;
wire  I_1644_D;
wire  I_1645_D;
wire  I_1645_G;
wire  I_1648_D;
wire  I_1649_D;
wire  I_1650_D;
wire  I_1651_D;
wire  I_1651_G;
wire  I_1660_D;
wire  I_1662_D;
wire  I_1667_D;
wire  I_1668_D;
wire  I_1671_S;
wire  I_1672_D;
wire  I_1673_D;
wire  I_1674_D;
wire  I_1674_S;
wire  I_1675_D;
wire  I_1675_G;
wire  I_1675_S;
wire  I_1676_D;
wire  I_1676_S;
wire  I_1677_D;
wire  I_1677_G;
wire  I_1677_S;
wire  I_1678_D;
wire  I_1679_D;
wire  I_1681_S;
wire  I_1682_D;
wire  I_1682_S;
wire  I_1683_D;
wire  I_1683_G;
wire  I_1683_S;
wire  I_1684_S;
wire  I_1685_D;
wire  I_1685_G;
wire  I_1685_S;
wire  I_1687_S;
wire  I_1689_D;
wire  I_168_D;
wire  I_1692_D;
wire  I_1693_D;
wire  I_1694_D;
wire  I_1695_D;
wire  I_1697_D;
wire  I_1699_D;
wire  I_169_D;
wire  I_169_G;
wire  I_16_D;
wire  I_1701_D;
wire  I_1706_D;
wire  I_1706_G;
wire  I_1707_D;
wire  I_1709_D;
wire  I_1713_D;
wire  I_1715_D;
wire  I_1729_D;
wire  I_1729_S;
wire  I_172_D;
wire  I_1730_G;
wire  I_1731_D;
wire  I_1731_S;
wire  I_1733_D;
wire  I_1733_S;
wire  I_1735_D;
wire  I_1735_S;
wire  I_1736_D;
wire  I_1737_D;
wire  I_1738_D;
wire  I_1738_G;
wire  I_1738_S;
wire  I_1739_D;
wire  I_1739_G;
wire  I_1739_S;
wire  I_173_D;
wire  I_173_G;
wire  I_1740_G;
wire  I_1740_S;
wire  I_1741_S;
wire  I_1742_D;
wire  I_1743_D;
wire  I_1744_G;
wire  I_1744_S;
wire  I_1746_G;
wire  I_1746_S;
wire  I_1748_S;
wire  I_1749_S;
wire  I_174_D;
wire  I_1750_S;
wire  I_1751_S;
wire  I_1752_S;
wire  I_1753_S;
wire  I_1755_D;
wire  I_1757_D;
wire  I_1758_S;
wire  I_1759_S;
wire  I_175_D;
wire  I_175_G;
wire  I_1761_D;
wire  I_1761_G;
wire  I_1763_D;
wire  I_176_D;
wire  I_1770_D;
wire  I_1771_D;
wire  I_1771_G;
wire  I_1772_D;
wire  I_1773_D;
wire  I_1773_G;
wire  I_1778_D;
wire  I_1779_D;
wire  I_1779_G;
wire  I_177_D;
wire  I_177_G;
wire  I_178_D;
wire  I_1798_D;
wire  I_179_D;
wire  I_179_G;
wire  I_17_D;
wire  I_17_G;
wire  I_1800_D;
wire  I_1802_D;
wire  I_1803_D;
wire  I_1803_G;
wire  I_1804_D;
wire  I_1805_D;
wire  I_1805_G;
wire  I_1806_D;
wire  I_1807_D;
wire  I_1808_D;
wire  I_1810_D;
wire  I_1811_D;
wire  I_1811_G;
wire  I_1812_D;
wire  I_1821_D;
wire  I_1822_D;
wire  I_1825_D;
wire  I_1826_D;
wire  I_1828_D;
wire  I_1831_S;
wire  I_1832_D;
wire  I_1832_S;
wire  I_1833_G;
wire  I_1833_S;
wire  I_1834_D;
wire  I_1834_S;
wire  I_1835_D;
wire  I_1835_G;
wire  I_1835_S;
wire  I_1836_D;
wire  I_1836_S;
wire  I_1837_D;
wire  I_1837_G;
wire  I_1837_S;
wire  I_1839_S;
wire  I_1843_S;
wire  I_1844_D;
wire  I_1845_D;
wire  I_1847_D;
wire  I_1853_S;
wire  I_1854_D;
wire  I_1855_D;
wire  I_1858_D;
wire  I_185_D;
wire  I_1861_D;
wire  I_1864_D;
wire  I_1864_G;
wire  I_1865_D;
wire  I_1870_D;
wire  I_1870_G;
wire  I_1871_D;
wire  I_1873_D;
wire  I_1874_D;
wire  I_1874_G;
wire  I_1876_D;
wire  I_1876_G;
wire  I_1879_D;
wire  I_1881_D;
wire  I_1888_D;
wire  I_1888_G;
wire  I_1889_D;
wire  I_1890_D;
wire  I_1891_S;
wire  I_1893_D;
wire  I_1893_S;
wire  I_1895_D;
wire  I_1895_S;
wire  I_1896_D;
wire  I_1896_G;
wire  I_1896_S;
wire  I_1897_D;
wire  I_1897_G;
wire  I_1897_S;
wire  I_1899_D;
wire  I_1899_S;
wire  I_18_D;
wire  I_1900_D;
wire  I_1901_D;
wire  I_1902_D;
wire  I_1902_G;
wire  I_1902_S;
wire  I_1903_D;
wire  I_1903_G;
wire  I_1903_S;
wire  I_1904_G;
wire  I_1904_S;
wire  I_1906_S;
wire  I_1907_G;
wire  I_1907_S;
wire  I_1908_S;
wire  I_1909_G;
wire  I_1909_S;
wire  I_190_D;
wire  I_1911_D;
wire  I_1911_S;
wire  I_1913_D;
wire  I_1913_S;
wire  I_1915_D;
wire  I_1915_S;
wire  I_1916_D;
wire  I_1917_D;
wire  I_1919_D;
wire  I_191_D;
wire  I_191_G;
wire  I_1921_G;
wire  I_1923_D;
wire  I_1928_D;
wire  I_1929_D;
wire  I_1929_G;
wire  I_1934_D;
wire  I_1935_D;
wire  I_1935_G;
wire  I_1936_D;
wire  I_1937_D;
wire  I_1937_G;
wire  I_1938_D;
wire  I_1939_D;
wire  I_1939_G;
wire  I_193_D;
wire  I_1943_D;
wire  I_1946_D;
wire  I_1947_D;
wire  I_1947_G;
wire  I_1949_D;
wire  I_1952_D;
wire  I_1958_D;
wire  I_1960_D;
wire  I_1961_D;
wire  I_1961_G;
wire  I_1962_D;
wire  I_1969_D;
wire  I_196_D;
wire  I_1970_D;
wire  I_1971_D;
wire  I_1971_G;
wire  I_1973_D;
wire  I_1982_D;
wire  I_1985_S;
wire  I_1986_D;
wire  I_1987_D;
wire  I_1988_D;
wire  I_1991_S;
wire  I_1992_D;
wire  I_1992_S;
wire  I_1993_D;
wire  I_1993_G;
wire  I_1993_S;
wire  I_1994_D;
wire  I_1995_S;
wire  I_1997_D;
wire  I_1998_D;
wire  I_1999_D;
wire  I_19_D;
wire  I_19_G;
wire  I_2001_S;
wire  I_2002_D;
wire  I_2002_S;
wire  I_2003_D;
wire  I_2003_G;
wire  I_2003_S;
wire  I_2004_S;
wire  I_2005_G;
wire  I_2005_S;
wire  I_2007_D;
wire  I_2009_D;
wire  I_200_D;
wire  I_2010_D;
wire  I_2011_D;
wire  I_2012_D;
wire  I_2013_D;
wire  I_2014_D;
wire  I_2015_D;
wire  I_201_D;
wire  I_201_G;
wire  I_2021_D;
wire  I_2024_D;
wire  I_2024_G;
wire  I_2025_D;
wire  I_2026_D;
wire  I_2026_G;
wire  I_2028_D;
wire  I_2028_G;
wire  I_2029_D;
wire  I_202_D;
wire  I_2033_D;
wire  I_2034_D;
wire  I_2034_G;
wire  I_2035_D;
wire  I_2041_D;
wire  I_2049_D;
wire  I_204_D;
wire  I_2050_D;
wire  I_2050_G;
wire  I_2051_D;
wire  I_2053_D;
wire  I_2053_S;
wire  I_2055_D;
wire  I_2055_S;
wire  I_2056_D;
wire  I_2056_G;
wire  I_2056_S;
wire  I_2057_D;
wire  I_2057_G;
wire  I_2057_S;
wire  I_2058_S;
wire  I_2059_G;
wire  I_2059_S;
wire  I_205_D;
wire  I_205_G;
wire  I_2060_D;
wire  I_2060_G;
wire  I_2060_S;
wire  I_2061_D;
wire  I_2061_G;
wire  I_2061_S;
wire  I_2062_D;
wire  I_2062_G;
wire  I_2063_D;
wire  I_2065_S;
wire  I_2066_D;
wire  I_2066_G;
wire  I_2066_S;
wire  I_2067_D;
wire  I_2067_G;
wire  I_2067_S;
wire  I_2068_D;
wire  I_2069_D;
wire  I_206_D;
wire  I_2071_D;
wire  I_2071_S;
wire  I_2073_D;
wire  I_2074_D;
wire  I_2075_D;
wire  I_2076_D;
wire  I_2077_D;
wire  I_2078_S;
wire  I_2079_S;
wire  I_207_D;
wire  I_207_G;
wire  I_2083_G;
wire  I_2088_D;
wire  I_2089_D;
wire  I_2089_G;
wire  I_208_D;
wire  I_2092_D;
wire  I_2093_D;
wire  I_2093_G;
wire  I_2096_D;
wire  I_2097_D;
wire  I_2097_G;
wire  I_2098_D;
wire  I_2099_D;
wire  I_2099_G;
wire  I_209_D;
wire  I_209_G;
wire  I_20_D;
wire  I_2103_D;
wire  I_2105_D;
wire  I_210_D;
wire  I_2112_D;
wire  I_2113_D;
wire  I_2113_G;
wire  I_2114_D;
wire  I_2115_D;
wire  I_2118_D;
wire  I_211_D;
wire  I_211_G;
wire  I_2120_D;
wire  I_2121_D;
wire  I_2121_G;
wire  I_2123_D;
wire  I_2124_D;
wire  I_2125_D;
wire  I_2125_G;
wire  I_2126_D;
wire  I_2127_D;
wire  I_2128_D;
wire  I_2129_D;
wire  I_2129_G;
wire  I_2130_D;
wire  I_2131_D;
wire  I_2131_G;
wire  I_2132_D;
wire  I_2133_D;
wire  I_2133_G;
wire  I_2135_G;
wire  I_2138_D;
wire  I_2139_D;
wire  I_2140_D;
wire  I_2142_D;
wire  I_2147_S;
wire  I_2148_D;
wire  I_2151_S;
wire  I_2152_D;
wire  I_2152_S;
wire  I_2153_D;
wire  I_2153_G;
wire  I_2153_S;
wire  I_2154_D;
wire  I_2155_D;
wire  I_2157_S;
wire  I_2159_S;
wire  I_2160_D;
wire  I_2160_S;
wire  I_2161_D;
wire  I_2161_G;
wire  I_2161_S;
wire  I_2162_D;
wire  I_2162_S;
wire  I_2163_D;
wire  I_2163_G;
wire  I_2163_S;
wire  I_2165_S;
wire  I_2167_S;
wire  I_2169_D;
wire  I_2171_S;
wire  I_2172_D;
wire  I_2173_D;
wire  I_2174_D;
wire  I_2175_D;
wire  I_2177_D;
wire  I_2181_D;
wire  I_2184_D;
wire  I_2184_G;
wire  I_2185_D;
wire  I_2187_D;
wire  I_2190_D;
wire  I_2190_G;
wire  I_2191_D;
wire  I_2194_D;
wire  I_2194_G;
wire  I_2195_D;
wire  I_2197_D;
wire  I_2199_D;
wire  I_21_D;
wire  I_21_G;
wire  I_2201_D;
wire  I_2209_D;
wire  I_2209_S;
wire  I_220_D;
wire  I_2210_D;
wire  I_2211_D;
wire  I_2213_D;
wire  I_2213_S;
wire  I_2215_D;
wire  I_2215_S;
wire  I_2216_D;
wire  I_2216_G;
wire  I_2216_S;
wire  I_2217_D;
wire  I_2217_G;
wire  I_2217_S;
wire  I_2218_G;
wire  I_2218_S;
wire  I_2219_S;
wire  I_2222_D;
wire  I_2222_G;
wire  I_2222_S;
wire  I_2223_D;
wire  I_2223_G;
wire  I_2223_S;
wire  I_2224_D;
wire  I_2225_D;
wire  I_2226_D;
wire  I_2226_G;
wire  I_2226_S;
wire  I_2227_D;
wire  I_2227_G;
wire  I_2227_S;
wire  I_2228_G;
wire  I_2228_S;
wire  I_222_D;
wire  I_2231_D;
wire  I_2231_S;
wire  I_2233_D;
wire  I_2234_D;
wire  I_2235_D;
wire  I_2236_D;
wire  I_2237_D;
wire  I_2238_S;
wire  I_2239_S;
wire  I_223_D;
wire  I_223_G;
wire  I_2241_G;
wire  I_2248_D;
wire  I_2249_D;
wire  I_2249_G;
wire  I_224_D;
wire  I_2253_D;
wire  I_2254_D;
wire  I_2255_D;
wire  I_2255_G;
wire  I_2258_D;
wire  I_2259_D;
wire  I_2259_G;
wire  I_225_D;
wire  I_2263_D;
wire  I_2265_D;
wire  I_2267_D;
wire  I_2269_D;
wire  I_226_D;
wire  I_2272_D;
wire  I_2274_D;
wire  I_2275_D;
wire  I_2278_D;
wire  I_227_D;
wire  I_2280_D;
wire  I_2281_D;
wire  I_2281_G;
wire  I_2282_D;
wire  I_2285_G;
wire  I_2288_D;
wire  I_2289_D;
wire  I_2290_D;
wire  I_2291_D;
wire  I_2291_G;
wire  I_2292_D;
wire  I_2295_G;
wire  I_229_S;
wire  I_2302_D;
wire  I_2305_S;
wire  I_2306_S;
wire  I_2307_G;
wire  I_2307_S;
wire  I_2308_D;
wire  I_230_D;
wire  I_2311_S;
wire  I_2312_D;
wire  I_2312_S;
wire  I_2313_D;
wire  I_2313_G;
wire  I_2313_S;
wire  I_2314_S;
wire  I_2315_G;
wire  I_2315_S;
wire  I_2317_S;
wire  I_2318_D;
wire  I_2319_D;
wire  I_2321_S;
wire  I_2322_D;
wire  I_2322_S;
wire  I_2323_D;
wire  I_2323_G;
wire  I_2323_S;
wire  I_2329_D;
wire  I_232_D;
wire  I_232_S;
wire  I_2330_D;
wire  I_2331_D;
wire  I_2332_D;
wire  I_2333_D;
wire  I_2334_D;
wire  I_2335_D;
wire  I_233_D;
wire  I_233_G;
wire  I_233_S;
wire  I_2341_D;
wire  I_2344_D;
wire  I_2344_G;
wire  I_2345_D;
wire  I_2348_D;
wire  I_2348_G;
wire  I_234_D;
wire  I_2353_D;
wire  I_2354_D;
wire  I_2354_G;
wire  I_2355_D;
wire  I_2357_D;
wire  I_235_D;
wire  I_2361_D;
wire  I_2369_D;
wire  I_236_D;
wire  I_236_S;
wire  I_2370_G;
wire  I_2371_D;
wire  I_2371_S;
wire  I_2373_D;
wire  I_2373_S;
wire  I_2375_D;
wire  I_2375_S;
wire  I_2376_D;
wire  I_2376_G;
wire  I_2376_S;
wire  I_2377_D;
wire  I_2377_G;
wire  I_2377_S;
wire  I_2379_D;
wire  I_2379_S;
wire  I_237_D;
wire  I_237_G;
wire  I_237_S;
wire  I_2381_G;
wire  I_2381_S;
wire  I_2382_D;
wire  I_2383_D;
wire  I_2384_G;
wire  I_2384_S;
wire  I_2386_D;
wire  I_2386_G;
wire  I_2386_S;
wire  I_2387_D;
wire  I_2387_G;
wire  I_2387_S;
wire  I_2388_G;
wire  I_2388_S;
wire  I_2389_S;
wire  I_238_D;
wire  I_238_S;
wire  I_2390_D;
wire  I_2391_D;
wire  I_2393_D;
wire  I_2394_D;
wire  I_2395_D;
wire  I_2396_D;
wire  I_2397_D;
wire  I_2399_D;
wire  I_239_D;
wire  I_239_G;
wire  I_239_S;
wire  I_23_G;
wire  I_2402_D;
wire  I_2403_D;
wire  I_2403_G;
wire  I_2408_D;
wire  I_2409_D;
wire  I_2409_G;
wire  I_240_D;
wire  I_240_S;
wire  I_2410_D;
wire  I_2411_D;
wire  I_2411_G;
wire  I_2412_D;
wire  I_2413_D;
wire  I_2413_G;
wire  I_2418_D;
wire  I_2419_D;
wire  I_2419_G;
wire  I_241_D;
wire  I_241_G;
wire  I_241_S;
wire  I_2420_D;
wire  I_2421_D;
wire  I_2421_G;
wire  I_2425_D;
wire  I_2427_D;
wire  I_2429_D;
wire  I_242_D;
wire  I_242_S;
wire  I_2432_D;
wire  I_2433_D;
wire  I_2433_G;
wire  I_2434_D;
wire  I_2435_D;
wire  I_2435_G;
wire  I_2438_D;
wire  I_243_D;
wire  I_243_G;
wire  I_243_S;
wire  I_2440_D;
wire  I_2441_D;
wire  I_2441_G;
wire  I_2442_D;
wire  I_2443_D;
wire  I_2443_G;
wire  I_2444_D;
wire  I_2445_D;
wire  I_2445_G;
wire  I_2446_D;
wire  I_2447_D;
wire  I_2448_D;
wire  I_2450_D;
wire  I_2451_D;
wire  I_2451_G;
wire  I_2453_D;
wire  I_2454_D;
wire  I_2455_D;
wire  I_245_D;
wire  I_2462_D;
wire  I_2466_D;
wire  I_2466_S;
wire  I_2467_D;
wire  I_2467_G;
wire  I_2467_S;
wire  I_2468_D;
wire  I_2471_S;
wire  I_2472_D;
wire  I_2472_S;
wire  I_2473_D;
wire  I_2473_G;
wire  I_2473_S;
wire  I_2474_D;
wire  I_2474_S;
wire  I_2475_D;
wire  I_2475_G;
wire  I_2475_S;
wire  I_2476_D;
wire  I_2476_S;
wire  I_2477_D;
wire  I_2477_G;
wire  I_2477_S;
wire  I_2479_S;
wire  I_247_D;
wire  I_2482_D;
wire  I_2482_S;
wire  I_2483_D;
wire  I_2483_G;
wire  I_2483_S;
wire  I_2485_S;
wire  I_2487_S;
wire  I_2489_D;
wire  I_2490_D;
wire  I_2491_D;
wire  I_2492_D;
wire  I_2493_D;
wire  I_2494_D;
wire  I_2495_D;
wire  I_2497_D;
wire  I_2498_D;
wire  I_2498_G;
wire  I_24_D;
wire  I_2501_D;
wire  I_2504_D;
wire  I_2504_G;
wire  I_2505_D;
wire  I_2509_D;
wire  I_2510_D;
wire  I_2510_G;
wire  I_2511_D;
wire  I_2513_D;
wire  I_2514_D;
wire  I_2514_G;
wire  I_2515_D;
wire  I_2517_D;
wire  I_2519_D;
wire  I_251_S;
wire  I_2521_D;
wire  I_2529_D;
wire  I_2529_S;
wire  I_2530_S;
wire  I_2531_G;
wire  I_2531_S;
wire  I_2533_D;
wire  I_2533_S;
wire  I_2534_G;
wire  I_2535_D;
wire  I_2535_G;
wire  I_2535_S;
wire  I_2536_D;
wire  I_2536_G;
wire  I_2536_S;
wire  I_2537_D;
wire  I_2537_G;
wire  I_2537_S;
wire  I_2539_D;
wire  I_2539_S;
wire  I_253_S;
wire  I_2540_G;
wire  I_2540_S;
wire  I_2542_D;
wire  I_2542_G;
wire  I_2542_S;
wire  I_2543_D;
wire  I_2543_G;
wire  I_2543_S;
wire  I_2544_G;
wire  I_2544_S;
wire  I_2545_S;
wire  I_2546_D;
wire  I_2546_G;
wire  I_2546_S;
wire  I_2547_D;
wire  I_2547_G;
wire  I_2547_S;
wire  I_2549_D;
wire  I_2549_S;
wire  I_254_D;
wire  I_254_S;
wire  I_2550_G;
wire  I_2550_S;
wire  I_2553_D;
wire  I_2554_D;
wire  I_2555_D;
wire  I_2556_D;
wire  I_2557_D;
wire  I_2558_S;
wire  I_2559_S;
wire  I_255_D;
wire  I_255_G;
wire  I_255_S;
wire  I_2561_G;
wire  I_2562_D;
wire  I_2563_D;
wire  I_2563_G;
wire  I_2572_D;
wire  I_2573_D;
wire  I_2573_G;
wire  I_2574_D;
wire  I_2575_D;
wire  I_2575_G;
wire  I_2576_D;
wire  I_2577_D;
wire  I_2577_G;
wire  I_2578_D;
wire  I_2579_D;
wire  I_2579_G;
wire  I_2580_D;
wire  I_2581_D;
wire  I_2581_G;
wire  I_2585_D;
wire  I_2592_D;
wire  I_2594_D;
wire  I_2595_D;
wire  I_2595_G;
wire  I_2598_D;
wire  I_25_D;
wire  I_25_G;
wire  I_2601_D;
wire  I_2603_D;
wire  I_2604_D;
wire  I_2605_D;
wire  I_2605_G;
wire  I_2606_D;
wire  I_2607_D;
wire  I_2607_G;
wire  I_2609_D;
wire  I_2610_D;
wire  I_2611_D;
wire  I_2611_G;
wire  I_2612_D;
wire  I_2613_D;
wire  I_2613_G;
wire  I_2614_D;
wire  I_2618_D;
wire  I_261_D;
wire  I_2620_D;
wire  I_2622_D;
wire  I_2625_S;
wire  I_2626_D;
wire  I_2626_S;
wire  I_2627_D;
wire  I_2627_G;
wire  I_2627_S;
wire  I_2628_D;
wire  I_2631_S;
wire  I_2632_D;
wire  I_2633_D;
wire  I_2634_D;
wire  I_2635_D;
wire  I_2636_D;
wire  I_2636_S;
wire  I_2637_D;
wire  I_2637_G;
wire  I_2637_S;
wire  I_2638_D;
wire  I_2638_S;
wire  I_2639_D;
wire  I_2639_G;
wire  I_2639_S;
wire  I_263_D;
wire  I_2641_S;
wire  I_2642_D;
wire  I_2642_S;
wire  I_2643_D;
wire  I_2643_G;
wire  I_2643_S;
wire  I_2644_D;
wire  I_2644_S;
wire  I_2645_D;
wire  I_2645_G;
wire  I_2645_S;
wire  I_2649_D;
wire  I_2650_D;
wire  I_2650_S;
wire  I_2651_G;
wire  I_2651_S;
wire  I_2652_D;
wire  I_2653_D;
wire  I_2654_D;
wire  I_2655_D;
wire  I_2657_D;
wire  I_2658_D;
wire  I_2658_G;
wire  I_2659_D;
wire  I_265_D;
wire  I_2661_D;
wire  I_2664_D;
wire  I_2664_G;
wire  I_2665_D;
wire  I_2668_D;
wire  I_2668_G;
wire  I_2669_D;
wire  I_266_D;
wire  I_266_G;
wire  I_2673_D;
wire  I_2674_D;
wire  I_2674_G;
wire  I_2675_D;
wire  I_2679_D;
wire  I_267_D;
wire  I_2681_D;
wire  I_2689_D;
wire  I_268_D;
wire  I_268_G;
wire  I_2690_D;
wire  I_2690_G;
wire  I_2690_S;
wire  I_2691_D;
wire  I_2691_G;
wire  I_2691_S;
wire  I_2693_D;
wire  I_2693_S;
wire  I_2695_D;
wire  I_2695_S;
wire  I_2696_D;
wire  I_2696_G;
wire  I_2696_S;
wire  I_2697_D;
wire  I_2697_G;
wire  I_2697_S;
wire  I_2698_D;
wire  I_2699_D;
wire  I_269_D;
wire  I_2700_D;
wire  I_2700_G;
wire  I_2700_S;
wire  I_2701_D;
wire  I_2701_G;
wire  I_2701_S;
wire  I_2705_S;
wire  I_2706_D;
wire  I_2706_G;
wire  I_2706_S;
wire  I_2707_D;
wire  I_2707_G;
wire  I_2707_S;
wire  I_2709_D;
wire  I_2709_S;
wire  I_270_D;
wire  I_270_G;
wire  I_2710_G;
wire  I_2710_S;
wire  I_2711_S;
wire  I_2713_D;
wire  I_2714_D;
wire  I_2715_D;
wire  I_2716_D;
wire  I_2717_D;
wire  I_2718_S;
wire  I_2719_S;
wire  I_271_D;
wire  I_2722_D;
wire  I_2723_D;
wire  I_2723_G;
wire  I_2728_D;
wire  I_2729_D;
wire  I_2729_G;
wire  I_272_D;
wire  I_272_G;
wire  I_2732_D;
wire  I_2733_D;
wire  I_2733_G;
wire  I_2735_D;
wire  I_2736_D;
wire  I_2737_D;
wire  I_2737_G;
wire  I_2738_D;
wire  I_2739_D;
wire  I_2739_G;
wire  I_273_D;
wire  I_2741_D;
wire  I_2742_D;
wire  I_2743_D;
wire  I_2743_G;
wire  I_2745_D;
wire  I_2747_D;
wire  I_2749_D;
wire  I_274_D;
wire  I_274_G;
wire  I_2752_D;
wire  I_2753_D;
wire  I_2753_G;
wire  I_2754_D;
wire  I_2755_D;
wire  I_2755_G;
wire  I_2758_D;
wire  I_275_D;
wire  I_2760_D;
wire  I_2761_D;
wire  I_2761_G;
wire  I_2763_D;
wire  I_2764_D;
wire  I_2765_D;
wire  I_2765_G;
wire  I_2767_G;
wire  I_2770_D;
wire  I_2771_D;
wire  I_2771_G;
wire  I_2773_G;
wire  I_2775_D;
wire  I_277_D;
wire  I_2782_D;
wire  I_2786_D;
wire  I_2786_S;
wire  I_2787_D;
wire  I_2787_G;
wire  I_2787_S;
wire  I_2788_D;
wire  I_2791_S;
wire  I_2792_D;
wire  I_2792_S;
wire  I_2793_D;
wire  I_2793_G;
wire  I_2793_S;
wire  I_2794_D;
wire  I_2795_D;
wire  I_2796_D;
wire  I_2796_S;
wire  I_2797_D;
wire  I_2797_G;
wire  I_2797_S;
wire  I_2799_S;
wire  I_279_D;
wire  I_2800_S;
wire  I_2801_G;
wire  I_2801_S;
wire  I_2805_S;
wire  I_2807_S;
wire  I_2809_D;
wire  I_2810_D;
wire  I_2811_D;
wire  I_2812_D;
wire  I_2813_D;
wire  I_2814_D;
wire  I_2815_D;
wire  I_2817_D;
wire  I_2818_D;
wire  I_2818_G;
wire  I_2819_D;
wire  I_281_D;
wire  I_2821_D;
wire  I_2824_D;
wire  I_2824_G;
wire  I_2825_D;
wire  I_2826_D;
wire  I_2826_G;
wire  I_2828_D;
wire  I_2828_G;
wire  I_2829_D;
wire  I_2830_D;
wire  I_2830_G;
wire  I_2831_D;
wire  I_2834_D;
wire  I_2834_G;
wire  I_2835_D;
wire  I_2837_D;
wire  I_2839_D;
wire  I_2841_D;
wire  I_2849_D;
wire  I_2849_S;
wire  I_2850_D;
wire  I_2850_G;
wire  I_2850_S;
wire  I_2851_D;
wire  I_2851_G;
wire  I_2851_S;
wire  I_2853_D;
wire  I_2853_S;
wire  I_2855_D;
wire  I_2855_S;
wire  I_2856_D;
wire  I_2856_G;
wire  I_2856_S;
wire  I_2857_D;
wire  I_2857_G;
wire  I_2857_S;
wire  I_2859_G;
wire  I_2859_S;
wire  I_285_D;
wire  I_2860_D;
wire  I_2860_G;
wire  I_2860_S;
wire  I_2861_D;
wire  I_2861_G;
wire  I_2861_S;
wire  I_2862_D;
wire  I_2862_G;
wire  I_2862_S;
wire  I_2863_D;
wire  I_2863_G;
wire  I_2863_S;
wire  I_2864_D;
wire  I_2865_D;
wire  I_2866_D;
wire  I_2866_G;
wire  I_2866_S;
wire  I_2867_D;
wire  I_2867_G;
wire  I_2867_S;
wire  I_2869_D;
wire  I_2871_D;
wire  I_2871_S;
wire  I_2873_D;
wire  I_2874_D;
wire  I_2875_D;
wire  I_2876_D;
wire  I_2877_D;
wire  I_2879_D;
wire  I_2881_G;
wire  I_2882_D;
wire  I_2883_D;
wire  I_2883_G;
wire  I_2889_D;
wire  I_288_D;
wire  I_2890_D;
wire  I_2893_D;
wire  I_2894_D;
wire  I_2895_D;
wire  I_2895_G;
wire  I_2898_D;
wire  I_2899_D;
wire  I_2899_G;
wire  I_289_D;
wire  I_2900_D;
wire  I_2901_D;
wire  I_2901_G;
wire  I_2902_D;
wire  I_2903_D;
wire  I_2903_G;
wire  I_2905_D;
wire  I_2907_D;
wire  I_290_D;
wire  I_2912_D;
wire  I_2914_D;
wire  I_2915_D;
wire  I_2915_G;
wire  I_2918_D;
wire  I_291_D;
wire  I_2922_D;
wire  I_2928_D;
wire  I_2929_D;
wire  I_2930_D;
wire  I_2931_D;
wire  I_2931_G;
wire  I_2932_D;
wire  I_2933_D;
wire  I_2933_G;
wire  I_2934_D;
wire  I_2935_D;
wire  I_2935_G;
wire  I_293_D;
wire  I_293_S;
wire  I_2940_D;
wire  I_2942_D;
wire  I_2945_S;
wire  I_2946_D;
wire  I_2946_S;
wire  I_2947_D;
wire  I_2947_G;
wire  I_2947_S;
wire  I_2948_D;
wire  I_2951_S;
wire  I_2952_D;
wire  I_2953_D;
wire  I_2954_D;
wire  I_2955_D;
wire  I_2956_D;
wire  I_2957_D;
wire  I_2958_S;
wire  I_2959_G;
wire  I_2959_S;
wire  I_295_D;
wire  I_2961_S;
wire  I_2962_D;
wire  I_2962_S;
wire  I_2963_D;
wire  I_2963_G;
wire  I_2963_S;
wire  I_2964_D;
wire  I_2964_S;
wire  I_2965_D;
wire  I_2965_G;
wire  I_2965_S;
wire  I_2966_D;
wire  I_2966_S;
wire  I_2967_D;
wire  I_2967_G;
wire  I_2967_S;
wire  I_2969_D;
wire  I_296_G;
wire  I_296_S;
wire  I_2970_D;
wire  I_2971_D;
wire  I_2972_D;
wire  I_2972_S;
wire  I_2973_G;
wire  I_2973_S;
wire  I_2974_D;
wire  I_2975_D;
wire  I_297_S;
wire  I_2981_D;
wire  I_2987_D;
wire  I_298_D;
wire  I_298_G;
wire  I_298_S;
wire  I_2993_D;
wire  I_299_D;
wire  I_299_G;
wire  I_299_S;
wire  I_3004_D;
wire  I_3004_G;
wire  I_3009_D;
wire  I_300_D;
wire  I_300_G;
wire  I_300_S;
wire  I_3010_D;
wire  I_3013_D;
wire  I_3013_S;
wire  I_3015_D;
wire  I_3015_S;
wire  I_3016_D;
wire  I_3017_D;
wire  I_3018_G;
wire  I_3018_S;
wire  I_3019_G;
wire  I_3019_S;
wire  I_301_D;
wire  I_301_G;
wire  I_301_S;
wire  I_3020_D;
wire  I_3021_D;
wire  I_3022_D;
wire  I_3023_D;
wire  I_3024_G;
wire  I_3024_S;
wire  I_3027_D;
wire  I_3029_D;
wire  I_302_D;
wire  I_302_G;
wire  I_302_S;
wire  I_3031_D;
wire  I_3031_S;
wire  I_3033_D;
wire  I_3034_D;
wire  I_3035_D;
wire  I_3036_G;
wire  I_3036_S;
wire  I_3037_G;
wire  I_3037_S;
wire  I_3038_S;
wire  I_3039_S;
wire  I_303_D;
wire  I_303_G;
wire  I_303_S;
wire  I_3042_D;
wire  I_304_D;
wire  I_304_G;
wire  I_304_S;
wire  I_3059_D;
wire  I_305_D;
wire  I_305_G;
wire  I_305_S;
wire  I_3061_D;
wire  I_3063_D;
wire  I_3065_D;
wire  I_306_D;
wire  I_306_G;
wire  I_306_S;
wire  I_3072_D;
wire  I_3073_D;
wire  I_3073_G;
wire  I_3074_D;
wire  I_3075_D;
wire  I_3078_D;
wire  I_307_D;
wire  I_307_G;
wire  I_307_S;
wire  I_3080_D;
wire  I_3082_D;
wire  I_3083_D;
wire  I_3084_D;
wire  I_3086_D;
wire  I_3087_D;
wire  I_3088_D;
wire  I_308_D;
wire  I_3091_G;
wire  I_3093_G;
wire  I_3095_G;
wire  I_3098_D;
wire  I_309_D;
wire  I_3100_D;
wire  I_3102_D;
wire  I_3106_S;
wire  I_3107_G;
wire  I_3107_S;
wire  I_3108_D;
wire  I_3111_S;
wire  I_3112_D;
wire  I_3112_S;
wire  I_3113_G;
wire  I_3113_S;
wire  I_3114_S;
wire  I_3115_G;
wire  I_3115_S;
wire  I_3116_D;
wire  I_3116_S;
wire  I_3117_G;
wire  I_3117_S;
wire  I_3119_S;
wire  I_311_D;
wire  I_3123_S;
wire  I_3125_S;
wire  I_3127_S;
wire  I_3129_D;
wire  I_3130_D;
wire  I_3130_S;
wire  I_3131_G;
wire  I_3131_S;
wire  I_3132_D;
wire  I_3133_D;
wire  I_3134_D;
wire  I_3135_D;
wire  I_3137_D;
wire  I_313_D;
wire  I_3141_D;
wire  I_3146_D;
wire  I_3146_G;
wire  I_3147_D;
wire  I_3148_D;
wire  I_3148_G;
wire  I_3149_D;
wire  I_3151_D;
wire  I_3153_D;
wire  I_3155_D;
wire  I_3157_D;
wire  I_3159_D;
wire  I_315_D;
wire  I_3163_D;
wire  I_3169_D;
wire  I_3169_S;
wire  I_3170_D;
wire  I_3171_D;
wire  I_3173_D;
wire  I_3173_S;
wire  I_3175_D;
wire  I_3175_S;
wire  I_3176_D;
wire  I_3177_D;
wire  I_3178_D;
wire  I_3178_G;
wire  I_3178_S;
wire  I_3179_D;
wire  I_3179_G;
wire  I_3179_S;
wire  I_317_D;
wire  I_3180_D;
wire  I_3180_S;
wire  I_3181_D;
wire  I_3181_G;
wire  I_3181_S;
wire  I_3182_G;
wire  I_3182_S;
wire  I_3184_G;
wire  I_3184_S;
wire  I_3185_S;
wire  I_3189_S;
wire  I_3191_D;
wire  I_3191_S;
wire  I_3192_D;
wire  I_3193_D;
wire  I_3194_G;
wire  I_3194_S;
wire  I_3195_G;
wire  I_3195_S;
wire  I_3196_D;
wire  I_3197_D;
wire  I_3198_S;
wire  I_3199_S;
wire  I_319_D;
wire  I_3201_G;
wire  I_3202_D;
wire  I_3203_D;
wire  I_3203_G;
wire  I_3210_D;
wire  I_3211_D;
wire  I_3211_G;
wire  I_3212_D;
wire  I_3213_D;
wire  I_3213_G;
wire  I_3216_D;
wire  I_3217_D;
wire  I_3217_G;
wire  I_3219_D;
wire  I_321_D;
wire  I_3220_D;
wire  I_3221_D;
wire  I_3221_G;
wire  I_3225_D;
wire  I_3229_D;
wire  I_3232_D;
wire  I_3234_D;
wire  I_3235_D;
wire  I_3235_G;
wire  I_3238_D;
wire  I_3241_D;
wire  I_3242_D;
wire  I_3243_D;
wire  I_3243_G;
wire  I_3244_D;
wire  I_3245_D;
wire  I_3245_G;
wire  I_3246_D;
wire  I_3249_D;
wire  I_3251_G;
wire  I_3254_D;
wire  I_3258_D;
wire  I_3262_D;
wire  I_3265_S;
wire  I_3266_D;
wire  I_3266_S;
wire  I_3267_D;
wire  I_3267_G;
wire  I_3267_S;
wire  I_3268_D;
wire  I_3271_S;
wire  I_3276_D;
wire  I_3276_S;
wire  I_3277_D;
wire  I_3277_G;
wire  I_3277_S;
wire  I_3281_S;
wire  I_3283_S;
wire  I_3284_D;
wire  I_3285_D;
wire  I_3286_D;
wire  I_3287_D;
wire  I_3288_D;
wire  I_3289_D;
wire  I_3290_D;
wire  I_3291_D;
wire  I_3292_D;
wire  I_3293_D;
wire  I_3294_D;
wire  I_3295_D;
wire  I_329_D;
wire  I_32_D;
wire  I_3301_D;
wire  I_3308_D;
wire  I_3308_G;
wire  I_3309_D;
wire  I_3311_D;
wire  I_3313_D;
wire  I_3329_D;
wire  I_332_D;
wire  I_3331_D;
wire  I_3331_G;
wire  I_3333_D;
wire  I_3333_S;
wire  I_3335_D;
wire  I_3335_S;
wire  I_3337_D;
wire  I_3339_D;
wire  I_333_D;
wire  I_333_G;
wire  I_3340_D;
wire  I_3340_G;
wire  I_3340_S;
wire  I_3341_D;
wire  I_3341_G;
wire  I_3341_S;
wire  I_3342_G;
wire  I_3342_S;
wire  I_3345_D;
wire  I_3345_S;
wire  I_3347_D;
wire  I_3348_D;
wire  I_3349_D;
wire  I_334_D;
wire  I_3350_S;
wire  I_3351_S;
wire  I_3352_D;
wire  I_3353_D;
wire  I_3354_S;
wire  I_3355_S;
wire  I_3356_D;
wire  I_3357_D;
wire  I_3359_D;
wire  I_335_D;
wire  I_335_G;
wire  I_3363_D;
wire  I_3369_D;
wire  I_336_D;
wire  I_3371_D;
wire  I_3374_D;
wire  I_3375_D;
wire  I_3375_G;
wire  I_3376_D;
wire  I_3377_D;
wire  I_3377_G;
wire  I_3379_D;
wire  I_337_D;
wire  I_337_G;
wire  I_3381_G;
wire  I_338_D;
wire  I_3392_D;
wire  I_3393_D;
wire  I_3393_G;
wire  I_3398_D;
wire  I_339_D;
wire  I_339_G;
wire  I_33_D;
wire  I_3401_G;
wire  I_3403_G;
wire  I_3407_D;
wire  I_3408_D;
wire  I_3409_D;
wire  I_3409_G;
wire  I_3411_G;
wire  I_3412_D;
wire  I_3413_D;
wire  I_3414_D;
wire  I_3416_D;
wire  I_3418_D;
wire  I_341_D;
wire  I_3420_D;
wire  I_3423_D;
wire  I_3426_D;
wire  I_3427_D;
wire  I_3428_D;
wire  I_3431_S;
wire  I_3433_S;
wire  I_3435_S;
wire  I_3436_D;
wire  I_3439_S;
wire  I_3440_D;
wire  I_3440_S;
wire  I_3441_D;
wire  I_3441_G;
wire  I_3441_S;
wire  I_3443_S;
wire  I_3445_S;
wire  I_3446_D;
wire  I_3447_D;
wire  I_3448_D;
wire  I_3449_D;
wire  I_3450_D;
wire  I_3451_D;
wire  I_3452_D;
wire  I_3453_D;
wire  I_3454_S;
wire  I_3455_G;
wire  I_3455_S;
wire  I_3457_D;
wire  I_3461_D;
wire  I_3465_D;
wire  I_3467_D;
wire  I_3471_D;
wire  I_3475_D;
wire  I_3476_D;
wire  I_3476_G;
wire  I_3477_D;
wire  I_347_D;
wire  I_3480_D;
wire  I_3480_G;
wire  I_3481_D;
wire  I_3489_D;
wire  I_3489_S;
wire  I_3491_D;
wire  I_3491_S;
wire  I_3493_D;
wire  I_3493_S;
wire  I_3495_D;
wire  I_3495_S;
wire  I_3497_S;
wire  I_3499_D;
wire  I_3499_S;
wire  I_3500_D;
wire  I_3501_D;
wire  I_3503_D;
wire  I_3503_S;
wire  I_3504_D;
wire  I_3505_D;
wire  I_3507_D;
wire  I_3508_D;
wire  I_3508_G;
wire  I_3508_S;
wire  I_3509_D;
wire  I_3509_G;
wire  I_3509_S;
wire  I_3510_S;
wire  I_3511_S;
wire  I_3512_D;
wire  I_3512_G;
wire  I_3512_S;
wire  I_3513_D;
wire  I_3513_G;
wire  I_3513_S;
wire  I_3514_S;
wire  I_3515_S;
wire  I_3516_D;
wire  I_3517_D;
wire  I_3519_D;
wire  I_3521_D;
wire  I_3529_D;
wire  I_3529_G;
wire  I_3535_D;
wire  I_3538_D;
wire  I_3539_D;
wire  I_3539_G;
wire  I_3540_D;
wire  I_3541_D;
wire  I_3541_G;
wire  I_3549_D;
wire  I_354_D;
wire  I_3554_D;
wire  I_3555_G;
wire  I_3558_D;
wire  I_355_D;
wire  I_3561_G;
wire  I_3562_D;
wire  I_3563_D;
wire  I_3564_D;
wire  I_3565_D;
wire  I_3567_G;
wire  I_3568_D;
wire  I_3569_D;
wire  I_356_D;
wire  I_3570_D;
wire  I_3571_D;
wire  I_3571_G;
wire  I_3572_D;
wire  I_3573_D;
wire  I_3573_G;
wire  I_3574_D;
wire  I_3576_D;
wire  I_3578_D;
wire  I_3582_D;
wire  I_3584_D;
wire  I_3585_D;
wire  I_3586_D;
wire  I_3587_D;
wire  I_3588_D;
wire  I_3591_S;
wire  I_3593_G;
wire  I_3593_S;
wire  I_3595_S;
wire  I_3597_S;
wire  I_3599_S;
wire  I_3601_S;
wire  I_3602_D;
wire  I_3602_S;
wire  I_3603_D;
wire  I_3603_G;
wire  I_3603_S;
wire  I_3604_D;
wire  I_3604_S;
wire  I_3605_D;
wire  I_3605_G;
wire  I_3605_S;
wire  I_3606_D;
wire  I_3607_D;
wire  I_3608_D;
wire  I_3609_D;
wire  I_3610_D;
wire  I_3611_D;
wire  I_3612_D;
wire  I_3613_D;
wire  I_3614_D;
wire  I_3615_D;
wire  I_361_G;
wire  I_3621_D;
wire  I_3627_D;
wire  I_362_D;
wire  I_3633_D;
wire  I_3638_D;
wire  I_3638_G;
wire  I_3639_D;
wire  I_3649_D;
wire  I_3649_G;
wire  I_364_D;
wire  I_3651_D;
wire  I_3653_D;
wire  I_3653_S;
wire  I_3655_D;
wire  I_3655_S;
wire  I_3657_D;
wire  I_3658_G;
wire  I_3658_S;
wire  I_3659_G;
wire  I_3659_S;
wire  I_365_D;
wire  I_365_G;
wire  I_3660_D;
wire  I_3663_D;
wire  I_3663_S;
wire  I_3664_G;
wire  I_3664_S;
wire  I_3667_D;
wire  I_3667_S;
wire  I_3669_D;
wire  I_3669_S;
wire  I_366_D;
wire  I_3670_D;
wire  I_3670_G;
wire  I_3670_S;
wire  I_3671_D;
wire  I_3671_G;
wire  I_3671_S;
wire  I_3672_S;
wire  I_3673_S;
wire  I_3675_D;
wire  I_3676_D;
wire  I_3677_D;
wire  I_3678_S;
wire  I_3679_S;
wire  I_367_D;
wire  I_367_G;
wire  I_3681_D;
wire  I_3683_D;
wire  I_368_D;
wire  I_3691_D;
wire  I_3692_D;
wire  I_3695_D;
wire  I_3699_D;
wire  I_369_D;
wire  I_369_G;
wire  I_36_D;
wire  I_3701_D;
wire  I_3703_D;
wire  I_370_D;
wire  I_3718_D;
wire  I_371_D;
wire  I_371_G;
wire  I_3720_D;
wire  I_3724_D;
wire  I_3725_D;
wire  I_3727_G;
wire  I_3728_D;
wire  I_372_D;
wire  I_3731_G;
wire  I_3733_G;
wire  I_3735_G;
wire  I_3736_D;
wire  I_3738_D;
wire  I_373_D;
wire  I_3740_D;
wire  I_3742_D;
wire  I_3744_D;
wire  I_3745_D;
wire  I_3746_D;
wire  I_3747_D;
wire  I_3748_D;
wire  I_3751_S;
wire  I_3752_D;
wire  I_3753_D;
wire  I_3755_D;
wire  I_3755_S;
wire  I_3759_S;
wire  I_375_D;
wire  I_3763_S;
wire  I_3765_S;
wire  I_3766_D;
wire  I_3767_D;
wire  I_3767_G;
wire  I_3768_D;
wire  I_3769_D;
wire  I_3770_D;
wire  I_3771_D;
wire  I_3772_D;
wire  I_3773_D;
wire  I_3774_D;
wire  I_3775_D;
wire  I_3781_D;
wire  I_3788_D;
wire  I_3791_D;
wire  I_3793_D;
wire  I_3795_D;
wire  I_3797_D;
wire  I_379_G;
wire  I_3808_D;
wire  I_3809_D;
wire  I_3810_D;
wire  I_3811_D;
wire  I_3813_D;
wire  I_3813_S;
wire  I_3815_D;
wire  I_3815_S;
wire  I_3816_D;
wire  I_3817_D;
wire  I_3818_D;
wire  I_3819_G;
wire  I_381_G;
wire  I_3820_D;
wire  I_3823_D;
wire  I_3823_S;
wire  I_3824_G;
wire  I_3824_S;
wire  I_3825_D;
wire  I_3825_S;
wire  I_3827_D;
wire  I_3829_D;
wire  I_3829_S;
wire  I_382_D;
wire  I_3830_D;
wire  I_3830_G;
wire  I_3831_D;
wire  I_3832_S;
wire  I_3833_S;
wire  I_3834_D;
wire  I_3835_D;
wire  I_3836_D;
wire  I_3836_G;
wire  I_3837_D;
wire  I_3838_S;
wire  I_3839_S;
wire  I_3845_D;
wire  I_3847_D;
wire  I_3847_G;
wire  I_3850_D;
wire  I_3851_G;
wire  I_3852_D;
wire  I_3854_D;
wire  I_3855_D;
wire  I_3855_G;
wire  I_3856_D;
wire  I_3857_D;
wire  I_3857_G;
wire  I_3859_D;
wire  I_385_D;
wire  I_3861_D;
wire  I_3867_D;
wire  I_3869_D;
wire  I_3872_D;
wire  I_3874_D;
wire  I_387_S;
wire  I_3880_D;
wire  I_3882_D;
wire  I_3883_D;
wire  I_3884_D;
wire  I_3887_D;
wire  I_3889_D;
wire  I_3893_G;
wire  I_3894_D;
wire  I_3896_D;
wire  I_389_S;
wire  I_3902_D;
wire  I_3904_D;
wire  I_3904_S;
wire  I_3905_G;
wire  I_3905_S;
wire  I_3906_D;
wire  I_3906_S;
wire  I_3907_G;
wire  I_3907_S;
wire  I_3908_D;
wire  I_3909_D;
wire  I_390_D;
wire  I_3910_D;
wire  I_3911_D;
wire  I_3911_G;
wire  I_3912_D;
wire  I_3913_S;
wire  I_3915_G;
wire  I_3915_S;
wire  I_3917_S;
wire  I_3919_S;
wire  I_3921_S;
wire  I_3923_G;
wire  I_3923_S;
wire  I_3924_D;
wire  I_3924_S;
wire  I_3925_D;
wire  I_3925_G;
wire  I_3925_S;
wire  I_3926_D;
wire  I_3926_S;
wire  I_3927_G;
wire  I_3927_S;
wire  I_3928_D;
wire  I_3929_D;
wire  I_3930_D;
wire  I_3931_D;
wire  I_3932_D;
wire  I_3933_D;
wire  I_3933_G;
wire  I_3934_D;
wire  I_3935_D;
wire  I_3937_D;
wire  I_3939_D;
wire  I_393_S;
wire  I_394_D;
wire  I_3950_D;
wire  I_3950_G;
wire  I_3953_D;
wire  I_3955_D;
wire  I_3956_D;
wire  I_3956_G;
wire  I_3958_D;
wire  I_3958_G;
wire  I_395_D;
wire  I_3961_D;
wire  I_3968_G;
wire  I_3968_S;
wire  I_3969_S;
wire  I_396_D;
wire  I_396_S;
wire  I_3970_G;
wire  I_3970_S;
wire  I_3971_G;
wire  I_3971_S;
wire  I_3972_D;
wire  I_3973_D;
wire  I_3974_D;
wire  I_3974_G;
wire  I_3975_D;
wire  I_3976_D;
wire  I_3977_D;
wire  I_3977_G;
wire  I_3979_D;
wire  I_397_D;
wire  I_397_G;
wire  I_397_S;
wire  I_3980_D;
wire  I_3980_G;
wire  I_3981_D;
wire  I_3982_G;
wire  I_3983_D;
wire  I_3983_G;
wire  I_3983_S;
wire  I_3985_D;
wire  I_3985_S;
wire  I_3986_G;
wire  I_3986_S;
wire  I_3987_G;
wire  I_3987_S;
wire  I_3988_G;
wire  I_3988_S;
wire  I_3989_G;
wire  I_3989_S;
wire  I_398_D;
wire  I_398_S;
wire  I_3990_G;
wire  I_3990_S;
wire  I_3991_G;
wire  I_3991_S;
wire  I_3992_G;
wire  I_3992_S;
wire  I_3993_G;
wire  I_3993_S;
wire  I_3994_D;
wire  I_3995_D;
wire  I_3996_D;
wire  I_3997_D;
wire  I_3999_D;
wire  I_3999_G;
wire  I_399_D;
wire  I_399_G;
wire  I_399_S;
wire  I_3_D;
wire  I_3_G;
wire  I_400_D;
wire  I_400_S;
wire  I_401_D;
wire  I_401_G;
wire  I_401_S;
wire  I_402_D;
wire  I_402_S;
wire  I_403_D;
wire  I_403_G;
wire  I_403_S;
wire  I_404_S;
wire  I_405_G;
wire  I_405_S;
wire  I_409_S;
wire  I_40_D;
wire  I_410_D;
wire  I_410_S;
wire  I_411_D;
wire  I_411_G;
wire  I_411_S;
wire  I_415_S;
wire  I_418_D;
wire  I_418_G;
wire  I_419_D;
wire  I_41_D;
wire  I_41_G;
wire  I_421_D;
wire  I_423_D;
wire  I_426_D;
wire  I_426_G;
wire  I_429_D;
wire  I_42_D;
wire  I_430_D;
wire  I_430_G;
wire  I_431_D;
wire  I_432_D;
wire  I_432_G;
wire  I_433_D;
wire  I_434_D;
wire  I_434_G;
wire  I_435_D;
wire  I_437_D;
wire  I_439_D;
wire  I_43_D;
wire  I_43_G;
wire  I_443_D;
wire  I_445_D;
wire  I_447_D;
wire  I_448_D;
wire  I_449_D;
wire  I_44_D;
wire  I_450_D;
wire  I_450_G;
wire  I_450_S;
wire  I_451_D;
wire  I_451_G;
wire  I_451_S;
wire  I_453_D;
wire  I_453_S;
wire  I_455_D;
wire  I_456_D;
wire  I_457_D;
wire  I_458_S;
wire  I_459_G;
wire  I_459_S;
wire  I_45_D;
wire  I_45_G;
wire  I_460_G;
wire  I_460_S;
wire  I_461_S;
wire  I_462_D;
wire  I_462_G;
wire  I_462_S;
wire  I_463_D;
wire  I_463_G;
wire  I_463_S;
wire  I_464_D;
wire  I_464_G;
wire  I_464_S;
wire  I_465_D;
wire  I_465_G;
wire  I_465_S;
wire  I_466_D;
wire  I_466_G;
wire  I_466_S;
wire  I_467_D;
wire  I_467_G;
wire  I_467_S;
wire  I_468_D;
wire  I_469_D;
wire  I_46_D;
wire  I_471_D;
wire  I_471_S;
wire  I_473_D;
wire  I_475_D;
wire  I_477_D;
wire  I_477_S;
wire  I_479_D;
wire  I_47_D;
wire  I_47_G;
wire  I_482_D;
wire  I_483_D;
wire  I_483_G;
wire  I_48_D;
wire  I_493_G;
wire  I_494_D;
wire  I_495_D;
wire  I_495_G;
wire  I_496_D;
wire  I_497_D;
wire  I_497_G;
wire  I_498_D;
wire  I_499_D;
wire  I_499_G;
wire  I_49_D;
wire  I_49_G;
wire  I_500_D;
wire  I_501_D;
wire  I_501_G;
wire  I_503_D;
wire  I_503_G;
wire  I_505_D;
wire  I_507_G;
wire  I_509_D;
wire  I_50_D;
wire  I_511_D;
wire  I_513_D;
wire  I_516_D;
wire  I_51_D;
wire  I_51_G;
wire  I_520_D;
wire  I_522_D;
wire  I_524_D;
wire  I_525_D;
wire  I_526_D;
wire  I_527_D;
wire  I_527_G;
wire  I_528_D;
wire  I_529_D;
wire  I_529_G;
wire  I_52_D;
wire  I_530_D;
wire  I_531_D;
wire  I_531_G;
wire  I_532_D;
wire  I_533_D;
wire  I_533_G;
wire  I_535_G;
wire  I_539_G;
wire  I_53_D;
wire  I_53_G;
wire  I_543_G;
wire  I_544_D;
wire  I_545_D;
wire  I_546_D;
wire  I_547_D;
wire  I_549_S;
wire  I_550_D;
wire  I_552_D;
wire  I_553_D;
wire  I_554_D;
wire  I_555_D;
wire  I_556_S;
wire  I_557_G;
wire  I_557_S;
wire  I_558_D;
wire  I_558_S;
wire  I_559_D;
wire  I_559_G;
wire  I_559_S;
wire  I_55_G;
wire  I_560_D;
wire  I_560_S;
wire  I_561_D;
wire  I_561_G;
wire  I_561_S;
wire  I_562_D;
wire  I_562_S;
wire  I_563_D;
wire  I_563_G;
wire  I_563_S;
wire  I_564_D;
wire  I_564_S;
wire  I_565_D;
wire  I_565_G;
wire  I_565_S;
wire  I_566_D;
wire  I_566_S;
wire  I_567_D;
wire  I_567_G;
wire  I_567_S;
wire  I_56_D;
wire  I_571_G;
wire  I_572_D;
wire  I_573_D;
wire  I_575_S;
wire  I_57_D;
wire  I_57_G;
wire  I_581_D;
wire  I_583_D;
wire  I_584_D;
wire  I_584_G;
wire  I_586_D;
wire  I_586_G;
wire  I_588_D;
wire  I_588_G;
wire  I_589_D;
wire  I_590_D;
wire  I_590_G;
wire  I_591_D;
wire  I_592_D;
wire  I_592_G;
wire  I_593_D;
wire  I_594_D;
wire  I_594_G;
wire  I_595_D;
wire  I_596_D;
wire  I_596_G;
wire  I_597_D;
wire  I_59_D;
wire  I_601_D;
wire  I_603_D;
wire  I_607_D;
wire  I_608_D;
wire  I_609_D;
wire  I_610_D;
wire  I_611_D;
wire  I_613_D;
wire  I_613_S;
wire  I_615_D;
wire  I_616_S;
wire  I_617_G;
wire  I_617_S;
wire  I_618_S;
wire  I_619_G;
wire  I_619_S;
wire  I_620_D;
wire  I_620_G;
wire  I_620_S;
wire  I_621_D;
wire  I_621_G;
wire  I_621_S;
wire  I_622_D;
wire  I_622_G;
wire  I_622_S;
wire  I_623_D;
wire  I_623_G;
wire  I_623_S;
wire  I_624_D;
wire  I_624_G;
wire  I_624_S;
wire  I_625_D;
wire  I_625_G;
wire  I_625_S;
wire  I_626_D;
wire  I_626_G;
wire  I_626_S;
wire  I_627_D;
wire  I_627_G;
wire  I_627_S;
wire  I_628_D;
wire  I_628_G;
wire  I_628_S;
wire  I_629_D;
wire  I_629_G;
wire  I_629_S;
wire  I_631_D;
wire  I_633_D;
wire  I_634_D;
wire  I_635_D;
wire  I_637_D;
wire  I_638_G;
wire  I_638_S;
wire  I_639_S;
wire  I_640_D;
wire  I_641_D;
wire  I_641_G;
wire  I_648_D;
wire  I_649_D;
wire  I_649_G;
wire  I_652_D;
wire  I_653_D;
wire  I_653_G;
wire  I_654_D;
wire  I_655_D;
wire  I_655_G;
wire  I_656_D;
wire  I_657_D;
wire  I_657_G;
wire  I_658_D;
wire  I_659_D;
wire  I_659_G;
wire  I_65_S;
wire  I_660_D;
wire  I_661_D;
wire  I_661_G;
wire  I_667_D;
wire  I_670_D;
wire  I_671_D;
wire  I_671_G;
wire  I_674_D;
wire  I_675_D;
wire  I_676_D;
wire  I_67_D;
wire  I_67_S;
wire  I_680_D;
wire  I_681_D;
wire  I_681_G;
wire  I_682_D;
wire  I_684_D;
wire  I_685_D;
wire  I_685_G;
wire  I_686_D;
wire  I_687_D;
wire  I_687_G;
wire  I_688_D;
wire  I_689_D;
wire  I_689_G;
wire  I_690_D;
wire  I_691_D;
wire  I_691_G;
wire  I_692_D;
wire  I_693_D;
wire  I_693_G;
wire  I_698_D;
wire  I_699_D;
wire  I_69_S;
wire  I_700_D;
wire  I_705_D;
wire  I_707_S;
wire  I_709_S;
wire  I_70_D;
wire  I_710_D;
wire  I_713_S;
wire  I_714_D;
wire  I_715_D;
wire  I_716_D;
wire  I_716_S;
wire  I_717_D;
wire  I_717_G;
wire  I_717_S;
wire  I_718_D;
wire  I_718_S;
wire  I_719_D;
wire  I_719_G;
wire  I_719_S;
wire  I_720_D;
wire  I_720_S;
wire  I_721_D;
wire  I_721_G;
wire  I_721_S;
wire  I_722_D;
wire  I_722_S;
wire  I_723_D;
wire  I_723_G;
wire  I_723_S;
wire  I_727_D;
wire  I_729_S;
wire  I_72_D;
wire  I_72_S;
wire  I_730_S;
wire  I_731_G;
wire  I_731_S;
wire  I_733_S;
wire  I_735_D;
wire  I_738_D;
wire  I_738_G;
wire  I_739_D;
wire  I_73_D;
wire  I_73_G;
wire  I_73_S;
wire  I_741_D;
wire  I_743_D;
wire  I_747_D;
wire  I_748_D;
wire  I_748_G;
wire  I_749_D;
wire  I_74_D;
wire  I_74_S;
wire  I_750_D;
wire  I_750_G;
wire  I_751_D;
wire  I_752_D;
wire  I_752_G;
wire  I_753_D;
wire  I_754_D;
wire  I_754_G;
wire  I_755_D;
wire  I_759_D;
wire  I_75_D;
wire  I_75_G;
wire  I_75_S;
wire  I_763_D;
wire  I_765_D;
wire  I_767_D;
wire  I_768_D;
wire  I_769_D;
wire  I_76_D;
wire  I_76_S;
wire  I_770_D;
wire  I_770_G;
wire  I_770_S;
wire  I_771_D;
wire  I_771_G;
wire  I_771_S;
wire  I_773_D;
wire  I_773_S;
wire  I_775_D;
wire  I_777_D;
wire  I_778_G;
wire  I_778_S;
wire  I_779_S;
wire  I_77_D;
wire  I_77_G;
wire  I_77_S;
wire  I_780_D;
wire  I_780_G;
wire  I_780_S;
wire  I_781_D;
wire  I_781_G;
wire  I_781_S;
wire  I_782_D;
wire  I_782_G;
wire  I_782_S;
wire  I_783_D;
wire  I_783_G;
wire  I_783_S;
wire  I_784_D;
wire  I_784_G;
wire  I_784_S;
wire  I_785_D;
wire  I_785_G;
wire  I_785_S;
wire  I_786_D;
wire  I_786_G;
wire  I_786_S;
wire  I_787_D;
wire  I_787_G;
wire  I_787_S;
wire  I_789_D;
wire  I_78_D;
wire  I_78_S;
wire  I_791_D;
wire  I_793_D;
wire  I_795_D;
wire  I_797_D;
wire  I_798_G;
wire  I_798_S;
wire  I_799_S;
wire  I_79_D;
wire  I_79_G;
wire  I_79_S;
wire  I_802_D;
wire  I_803_D;
wire  I_803_G;
wire  I_809_D;
wire  I_80_D;
wire  I_80_S;
wire  I_810_D;
wire  I_811_D;
wire  I_811_G;
wire  I_812_D;
wire  I_813_D;
wire  I_813_G;
wire  I_814_D;
wire  I_815_D;
wire  I_815_G;
wire  I_816_D;
wire  I_817_D;
wire  I_817_G;
wire  I_818_D;
wire  I_819_D;
wire  I_819_G;
wire  I_81_D;
wire  I_81_G;
wire  I_81_S;
wire  I_821_D;
wire  I_825_D;
wire  I_827_D;
wire  I_82_D;
wire  I_82_S;
wire  I_833_D;
wire  I_836_D;
wire  I_83_D;
wire  I_83_G;
wire  I_83_S;
wire  I_842_D;
wire  I_843_D;
wire  I_843_G;
wire  I_844_D;
wire  I_845_D;
wire  I_845_G;
wire  I_846_D;
wire  I_847_D;
wire  I_847_G;
wire  I_848_D;
wire  I_849_D;
wire  I_849_G;
wire  I_850_D;
wire  I_851_D;
wire  I_851_G;
wire  I_852_D;
wire  I_853_D;
wire  I_855_D;
wire  I_858_D;
wire  I_859_D;
wire  I_85_G;
wire  I_861_G;
wire  I_862_D;
wire  I_864_D;
wire  I_865_D;
wire  I_866_D;
wire  I_867_D;
wire  I_869_S;
wire  I_870_D;
wire  I_873_D;
wire  I_874_D;
wire  I_874_S;
wire  I_875_D;
wire  I_875_G;
wire  I_875_S;
wire  I_876_D;
wire  I_876_S;
wire  I_877_D;
wire  I_877_G;
wire  I_877_S;
wire  I_878_D;
wire  I_878_S;
wire  I_879_D;
wire  I_879_G;
wire  I_879_S;
wire  I_87_G;
wire  I_880_D;
wire  I_880_S;
wire  I_881_D;
wire  I_881_G;
wire  I_881_S;
wire  I_882_D;
wire  I_882_S;
wire  I_883_D;
wire  I_883_G;
wire  I_883_S;
wire  I_884_S;
wire  I_885_G;
wire  I_885_S;
wire  I_88_D;
wire  I_88_S;
wire  I_890_S;
wire  I_891_G;
wire  I_891_S;
wire  I_894_D;
wire  I_89_D;
wire  I_89_G;
wire  I_89_S;
wire  I_8_D;
wire  I_901_D;
wire  I_903_D;
wire  I_906_D;
wire  I_906_G;
wire  I_907_D;
wire  I_908_D;
wire  I_908_G;
wire  I_909_D;
wire  I_910_D;
wire  I_910_G;
wire  I_911_D;
wire  I_912_D;
wire  I_912_G;
wire  I_913_D;
wire  I_914_D;
wire  I_914_G;
wire  I_915_D;
wire  I_917_D;
wire  I_919_D;
wire  I_91_G;
wire  I_921_D;
wire  I_923_D;
wire  I_925_D;
wire  I_928_D;
wire  I_929_D;
wire  I_930_D;
wire  I_931_D;
wire  I_933_D;
wire  I_933_S;
wire  I_935_D;
wire  I_937_D;
wire  I_938_D;
wire  I_938_G;
wire  I_938_S;
wire  I_939_D;
wire  I_939_G;
wire  I_939_S;
wire  I_93_S;
wire  I_940_D;
wire  I_940_G;
wire  I_940_S;
wire  I_941_D;
wire  I_941_G;
wire  I_941_S;
wire  I_942_D;
wire  I_942_G;
wire  I_942_S;
wire  I_943_D;
wire  I_943_G;
wire  I_943_S;
wire  I_944_D;
wire  I_944_G;
wire  I_944_S;
wire  I_945_D;
wire  I_945_G;
wire  I_945_S;
wire  I_946_D;
wire  I_946_G;
wire  I_946_S;
wire  I_947_D;
wire  I_947_G;
wire  I_947_S;
wire  I_948_D;
wire  I_949_D;
wire  I_951_D;
wire  I_953_D;
wire  I_954_D;
wire  I_955_D;
wire  I_957_D;
wire  I_957_S;
wire  I_959_D;
wire  I_95_D;
wire  I_95_G;
wire  I_960_D;
wire  I_961_D;
wire  I_961_G;
wire  I_969_D;
wire  I_970_D;
wire  I_971_D;
wire  I_971_G;
wire  I_972_D;
wire  I_973_D;
wire  I_973_G;
wire  I_975_D;
wire  I_976_D;
wire  I_977_D;
wire  I_977_G;
wire  I_978_D;
wire  I_979_D;
wire  I_979_G;
wire  I_983_D;
wire  I_989_D;
wire  I_994_D;
wire  I_995_D;
wire  I_998_D;
wire  I_99_D;
wire  I_9_D;
wire  I_9_G;

  //--------------------------------------------------------------------------
  // Input assignments
  //--------------------------------------------------------------------------

  // Clock input drivers
  assign I_151_G = CLK;
  assign I_95_G  = !CLK;
  assign I_503_G = CLK;

  // Inverting input pin drivers
  assign I_3988_G = !A8;
  assign I_3990_G = !A9;
  assign I_3987_G = !A10;
  assign I_3195_G = !A11;
  assign I_3923_G = !A12;
  assign I_3593_G = !A13;
  assign I_3659_G = !A14;
  assign I_3982_G = !A15;
  assign I_91_G   = !D0;
  assign I_507_G  = !D1;
  assign I_87_G   = !D2;
  assign I_23_G   = !D3;
  assign I_85_G   = !D4;
  assign I_571_G  = !D5;
  assign I_3993_G = !D6;
  assign I_1260_G = !D7;
  assign I_3529_G = !RnW;
  assign I_3971_G = !nMAP;

  // Input from a non bonded pad, set to assumed passive value
  assign I_1313_G = VDD;

  // Tying this unconnected net low avoids a hang where SYNC resets the
  // CLK divider so that no further progress is possible.
  assign I_1408_G = VSS;

  //--------------------------------------------------------------------------
  // Netlist repairs
  //--------------------------------------------------------------------------

  // Repairing nets based on comments in 006_mjb_sorted.v
  assign I_3331_G = I_3884_D;
  assign I_3977_G = I_3971_S;
  assign I_3_G    = I_1025_D;
  assign I_1025_G = I_1889_D;
  assign I_1409_G = I_1889_D;
  assign I_1153_G = I_2371_S;
  assign I_1185_G = I_2275_D;
  assign I_1729_S = I_2275_D;
  assign I_493_G  = I_1185_D;
  assign I_1262_G = I_3585_D;
  assign I_1888_G = I_1507_D;
  assign I_2535_G = I_1507_D;
  assign I_3649_G = I_261_D;
  assign I_1730_G = I_245_D;
  assign I_1761_G = I_245_D;
  assign I_1258_G = I_245_D;
  assign I_1921_G = I_1825_D;
  assign I_2113_G = I_1825_D;
  assign I_2241_G = I_1825_D;
  assign I_2433_G = I_1825_D;
  assign I_2561_G = I_1825_D;
  assign I_2753_G = I_1825_D;
  assign I_2881_G = I_1825_D;
  assign I_3073_G = I_1825_D;
  assign I_3201_G = I_1825_D;
  assign I_3393_G = I_1825_D;
  assign I_3830_G = I_1671_S;
  assign I_2050_G = I_3075_D;
  assign I_2849_S = I_2657_D;
  assign I_3911_G = I_2471_S;
  assign I_2083_G = I_3363_D;
  assign I_3555_G = I_3657_D;
  assign I_2370_G = I_3657_D;
  assign I_1415_S = I_2489_D;
  assign I_1250_G = I_247_D;
  assign I_1311_G = I_1283_D;
  assign I_3999_G = I_3353_D;
  assign I_3836_G = I_1511_S;
  assign I_3036_G = I_3829_S;
  assign I_3933_G = I_3973_D;
  assign I_3735_G = I_1755_D;
  assign I_3915_G = I_3133_D;
  assign I_3980_G = I_1821_D;
  assign I_3974_G = I_1821_D;
  assign I_3851_G = I_3990_S;
  assign I_2231_D = I_1991_S;
  assign I_3767_G = I_3904_D;
  assign I_3667_S = I_3663_D;
  assign I_3819_G = I_3861_D;
  assign I_3847_G = I_3453_D;
  assign I_3381_G = I_3906_D;
  assign I_1631_G = I_3195_S;
  assign I_1235_D = I_1139_D;
  assign I_1193_G = I_1257_D;
  assign I_3019_G = I_2379_S;
  assign I_2534_G = I_2530_S;
  assign I_471_S  = I_631_D;
  assign I_2133_G = I_2151_S;
  assign I_2062_G = I_2791_S;

  //--------------------------------------------------------------------------

  generic_nmos I_0(.D(I_33_D), .G(I_3_G), .S(I_32_D));
  generic_pmos I_1(.D(VDD), .G(I_3_G), .S(I_33_D));
  generic_nmos I_10(.D(I_10_D), .G(I_11_G), .S(I_42_D));
  generic_nmos I_100(.D(I_101_D), .G(I_329_D), .S(I_133_D));
  generic_nmos I_1000(.D(VSS), .G(I_969_D), .S(I_1033_D));
  generic_pmos I_1001(.D(VDD), .G(I_969_D), .S(I_1033_D));
  generic_nmos I_1002(.D(I_1002_D), .G(I_1003_G), .S(I_1034_D));
  generic_pmos I_1003(.D(I_1003_D), .G(I_1003_G), .S(I_1035_D));
  generic_nmos I_1004(.D(I_1004_D), .G(I_1005_G), .S(I_1036_D));
  generic_pmos I_1005(.D(I_1005_D), .G(I_1005_G), .S(I_1037_D));
  generic_nmos I_1006(.D(VSS), .G(I_1997_D), .S(I_1038_D));
  generic_pmos I_1007(.D(VDD), .G(I_1997_D), .S(I_1039_D));
  generic_nmos I_1008(.D(I_1008_D), .G(I_1009_G), .S(I_1040_D));
  generic_pmos I_1009(.D(I_1009_D), .G(I_1009_G), .S(I_1041_D));
  generic_pmos I_101(.D(I_101_D), .G(I_395_D), .S(I_133_D));
  generic_nmos I_1010(.D(I_1010_D), .G(I_1011_G), .S(I_1042_D));
  generic_pmos I_1011(.D(I_1011_D), .G(I_1011_G), .S(I_1043_D));
  generic_nmos I_1012(.D(VSS), .G(I_983_D), .S(I_1045_D));
  generic_pmos I_1013(.D(VDD), .G(I_983_D), .S(I_1045_D));
  generic_nmos I_1014(.D(I_1014_D), .G(I_1113_S), .S(VSS));
  generic_pmos I_1015(.D(I_1015_D), .G(I_1113_S), .S(VDD));
  generic_nmos I_1016(.D(I_1401_D), .G(I_953_D), .S(VSS));
  generic_pmos I_1017(.D(I_1401_D), .G(I_953_D), .S(VDD));
  generic_nmos I_1018(.D(VSS), .G(I_1019_G), .S(VSS));
  generic_pmos I_1019(.D(VDD), .G(I_1019_G), .S(VDD));
  generic_nmos I_102(.D(I_103_D), .G(I_395_D), .S(I_135_D));
  generic_nmos I_1020(.D(VSS), .G(I_925_D), .S(I_1397_D));
  generic_pmos I_1021(.D(VDD), .G(I_925_D), .S(I_1397_D));
  generic_nmos I_1022(.D(I_1022_D), .G(I_1117_D), .S(VSS));
  generic_pmos I_1023(.D(I_1087_D), .G(I_1117_D), .S(VDD));
  generic_nmos I_1024(.D(I_1025_D), .G(I_1025_G), .S(VSS));
  generic_pmos I_1025(.D(I_1025_D), .G(I_1025_G), .S(VDD));
  generic_nmos I_1026(.D(VSS), .G(I_1249_D), .S(I_1027_S));
  generic_pmos I_1027(.D(VDD), .G(I_1249_D), .S(I_1027_S));
  generic_nmos I_1028(.D(I_1028_D), .G(I_1093_D), .S(I_1029_D));
  generic_pmos I_1029(.D(I_1029_D), .G(I_1093_D), .S(VDD));
  generic_pmos I_103(.D(I_103_D), .G(I_329_D), .S(I_135_D));
  generic_nmos I_1030(.D(VSS), .G(I_1095_D), .S(I_1093_S));
  generic_pmos I_1031(.D(VDD), .G(I_1095_D), .S(I_1093_S));
  generic_nmos I_1032(.D(I_1033_D), .G(I_969_D), .S(VSS));
  generic_pmos I_1033(.D(I_1033_D), .G(I_969_D), .S(VDD));
  generic_nmos I_1034(.D(I_1034_D), .G(I_1035_G), .S(I_1034_S));
  generic_pmos I_1035(.D(I_1035_D), .G(I_1035_G), .S(I_1035_S));
  generic_nmos I_1036(.D(I_1036_D), .G(I_1037_G), .S(I_1036_S));
  generic_pmos I_1037(.D(I_1037_D), .G(I_1037_G), .S(I_1037_S));
  generic_nmos I_1038(.D(I_1038_D), .G(I_1741_S), .S(I_1039_D));
  generic_pmos I_1039(.D(I_1039_D), .G(I_1741_S), .S(VDD));
  generic_nmos I_104(.D(I_104_D), .G(I_104_G), .S(I_136_D));
  generic_nmos I_1040(.D(I_1040_D), .G(I_1041_G), .S(I_1040_S));
  generic_pmos I_1041(.D(I_1041_D), .G(I_1041_G), .S(I_1041_S));
  generic_nmos I_1042(.D(I_1042_D), .G(I_1043_G), .S(I_1042_S));
  generic_pmos I_1043(.D(I_1043_D), .G(I_1043_G), .S(I_1043_S));
  generic_nmos I_1044(.D(I_1045_D), .G(I_983_D), .S(VSS));
  generic_pmos I_1045(.D(I_1045_D), .G(I_983_D), .S(VDD));
  generic_nmos I_1046(.D(VSS), .G(I_1047_G), .S(I_1046_S));
  generic_pmos I_1047(.D(VDD), .G(I_1047_G), .S(I_1047_S));
  generic_nmos I_1048(.D(VSS), .G(I_1401_D), .S(I_1049_S));
  generic_pmos I_1049(.D(VDD), .G(I_1401_D), .S(I_1049_S));
  generic_pmos I_105(.D(I_105_D), .G(I_136_G), .S(I_137_D));
  generic_nmos I_1050(.D(VSS), .G(I_445_D), .S(I_1051_S));
  generic_pmos I_1051(.D(VDD), .G(I_445_D), .S(I_1051_S));
  generic_nmos I_1052(.D(I_1397_D), .G(I_925_D), .S(VSS));
  generic_pmos I_1053(.D(I_1397_D), .G(I_925_D), .S(VDD));
  generic_nmos I_1054(.D(VSS), .G(I_1087_D), .S(I_1055_S));
  generic_pmos I_1055(.D(VDD), .G(I_1087_D), .S(I_1055_S));
  generic_nmos I_1056(.D(I_1089_D), .G(I_1153_G), .S(I_1088_D));
  generic_pmos I_1057(.D(VDD), .G(I_1667_D), .S(I_1089_D));
  generic_nmos I_1058(.D(I_1091_D), .G(I_389_S), .S(I_1090_D));
  generic_pmos I_1059(.D(VDD), .G(I_1985_S), .S(I_1091_D));
  generic_nmos I_106(.D(I_106_D), .G(I_106_G), .S(I_138_D));
  generic_nmos I_1060(.D(I_1061_D), .G(I_1097_S), .S(I_1093_D));
  generic_pmos I_1061(.D(I_1061_D), .G(I_715_D), .S(I_1093_D));
  generic_nmos I_1062(.D(I_1063_D), .G(I_715_D), .S(I_1095_D));
  generic_pmos I_1063(.D(I_1063_D), .G(I_1097_S), .S(I_1095_D));
  generic_nmos I_1064(.D(I_1097_S), .G(I_715_D), .S(VSS));
  generic_pmos I_1065(.D(I_1065_D), .G(I_1096_G), .S(VDD));
  generic_nmos I_1066(.D(I_1099_S), .G(I_1258_G), .S(VSS));
  generic_pmos I_1067(.D(I_1067_D), .G(I_1098_G), .S(VDD));
  generic_nmos I_1068(.D(I_1101_S), .G(I_1973_D), .S(VSS));
  generic_pmos I_1069(.D(I_1069_D), .G(I_1100_G), .S(VDD));
  generic_pmos I_107(.D(I_107_D), .G(I_138_G), .S(I_139_D));
  generic_nmos I_1070(.D(VSS), .G(I_975_D), .S(I_1102_D));
  generic_pmos I_1071(.D(VDD), .G(I_2471_S), .S(I_1103_D));
  generic_nmos I_1072(.D(I_1072_D), .G(I_1072_G), .S(I_1104_D));
  generic_pmos I_1073(.D(I_1073_D), .G(I_1104_G), .S(I_1105_D));
  generic_nmos I_1074(.D(I_1074_D), .G(I_1074_G), .S(I_1106_D));
  generic_pmos I_1075(.D(I_1075_D), .G(I_1106_G), .S(I_1107_D));
  generic_nmos I_1076(.D(I_1076_D), .G(I_1076_G), .S(I_1108_D));
  generic_pmos I_1077(.D(I_1077_D), .G(I_1108_G), .S(I_1109_D));
  generic_nmos I_1078(.D(I_2681_D), .G(I_1045_D), .S(I_1111_D));
  generic_pmos I_1079(.D(I_2681_D), .G(I_789_D), .S(I_1111_D));
  generic_nmos I_108(.D(I_108_D), .G(I_108_G), .S(I_140_D));
  generic_nmos I_1080(.D(VSS), .G(I_1529_D), .S(I_1112_D));
  generic_pmos I_1081(.D(VDD), .G(I_1529_D), .S(I_1113_D));
  generic_nmos I_1082(.D(I_1115_D), .G(I_1275_D), .S(I_1114_D));
  generic_pmos I_1083(.D(VDD), .G(I_1205_D), .S(I_1115_D));
  generic_nmos I_1084(.D(I_1117_D), .G(I_93_S), .S(I_1407_D));
  generic_pmos I_1085(.D(I_1085_D), .G(I_1116_G), .S(I_1117_D));
  generic_nmos I_1086(.D(I_1087_D), .G(I_95_D), .S(I_1119_D));
  generic_pmos I_1087(.D(I_1087_D), .G(I_93_S), .S(I_1119_D));
  generic_nmos I_1088(.D(I_1088_D), .G(I_1667_D), .S(VSS));
  generic_pmos I_1089(.D(I_1089_D), .G(I_1153_G), .S(VDD));
  generic_pmos I_109(.D(I_109_D), .G(I_140_G), .S(I_141_D));
  generic_nmos I_1090(.D(I_1090_D), .G(I_1985_S), .S(VSS));
  generic_pmos I_1091(.D(I_1091_D), .G(I_389_S), .S(VDD));
  generic_nmos I_1092(.D(I_1093_D), .G(I_715_D), .S(I_1093_S));
  generic_pmos I_1093(.D(I_1093_D), .G(I_1097_S), .S(I_1093_S));
  generic_nmos I_1094(.D(I_1095_D), .G(I_1097_S), .S(I_2169_D));
  generic_pmos I_1095(.D(I_1095_D), .G(I_715_D), .S(I_2169_D));
  generic_nmos I_1096(.D(VSS), .G(I_1096_G), .S(I_1096_S));
  generic_pmos I_1097(.D(VDD), .G(I_715_D), .S(I_1097_S));
  generic_nmos I_1098(.D(VSS), .G(I_1098_G), .S(I_1098_S));
  generic_pmos I_1099(.D(VDD), .G(I_1258_G), .S(I_1099_S));
  generic_pmos I_11(.D(I_11_D), .G(I_11_G), .S(I_43_D));
  generic_nmos I_110(.D(I_110_D), .G(I_110_G), .S(I_142_D));
  generic_nmos I_1100(.D(VSS), .G(I_1100_G), .S(I_1100_S));
  generic_pmos I_1101(.D(VDD), .G(I_1973_D), .S(I_1101_S));
  generic_nmos I_1102(.D(I_1102_D), .G(I_2471_S), .S(I_1103_D));
  generic_pmos I_1103(.D(I_1103_D), .G(I_975_D), .S(VDD));
  generic_nmos I_1104(.D(I_1104_D), .G(I_1104_G), .S(I_1104_S));
  generic_pmos I_1105(.D(I_1105_D), .G(I_1105_G), .S(I_1105_S));
  generic_nmos I_1106(.D(I_1106_D), .G(I_1106_G), .S(I_1106_S));
  generic_pmos I_1107(.D(I_1107_D), .G(I_1107_G), .S(I_1107_S));
  generic_nmos I_1108(.D(I_1108_D), .G(I_1108_G), .S(I_1108_S));
  generic_pmos I_1109(.D(I_1109_D), .G(I_1109_G), .S(I_1109_S));
  generic_pmos I_111(.D(I_111_D), .G(I_142_G), .S(I_143_D));
  generic_nmos I_1110(.D(I_1111_D), .G(I_789_D), .S(I_1207_D));
  generic_pmos I_1111(.D(I_1111_D), .G(I_1045_D), .S(I_1207_D));
  generic_nmos I_1112(.D(I_1112_D), .G(I_1529_D), .S(I_1113_S));
  generic_pmos I_1113(.D(I_1113_D), .G(I_1529_D), .S(I_1113_S));
  generic_nmos I_1114(.D(I_1114_D), .G(I_1205_D), .S(VSS));
  generic_pmos I_1115(.D(I_1115_D), .G(I_1275_D), .S(VDD));
  generic_nmos I_1116(.D(I_1407_D), .G(I_1116_G), .S(I_1116_S));
  generic_pmos I_1117(.D(I_1117_D), .G(I_95_D), .S(I_1407_D));
  generic_nmos I_1118(.D(I_1119_D), .G(I_93_S), .S(I_1247_D));
  generic_pmos I_1119(.D(I_1119_D), .G(I_95_D), .S(I_1247_D));
  generic_nmos I_112(.D(I_112_D), .G(I_112_G), .S(I_144_D));
  generic_nmos I_1120(.D(I_1120_D), .G(I_1121_G), .S(VSS));
  generic_pmos I_1121(.D(I_1121_D), .G(I_1121_G), .S(VDD));
  generic_nmos I_1122(.D(VSS), .G(I_1539_D), .S(I_1187_S));
  generic_pmos I_1123(.D(VDD), .G(I_1539_D), .S(I_1187_S));
  generic_nmos I_1124(.D(I_1221_D), .G(I_1189_D), .S(VSS));
  generic_pmos I_1125(.D(I_1221_D), .G(I_1189_D), .S(VDD));
  generic_nmos I_1126(.D(I_1223_D), .G(I_1187_S), .S(I_1158_D));
  generic_pmos I_1127(.D(VDD), .G(I_1187_S), .S(I_1223_D));
  generic_nmos I_1128(.D(I_1225_D), .G(I_1259_S), .S(VSS));
  generic_pmos I_1129(.D(I_1225_D), .G(I_1259_S), .S(VDD));
  generic_pmos I_113(.D(I_113_D), .G(I_144_G), .S(I_145_D));
  generic_nmos I_1130(.D(I_1227_D), .G(I_1195_D), .S(VSS));
  generic_pmos I_1131(.D(I_1227_D), .G(I_1195_D), .S(VDD));
  generic_nmos I_1132(.D(I_1132_D), .G(I_1133_G), .S(I_1164_D));
  generic_pmos I_1133(.D(I_1133_D), .G(I_1133_G), .S(I_1165_D));
  generic_nmos I_1134(.D(VSS), .G(I_1039_D), .S(I_1166_D));
  generic_pmos I_1135(.D(VDD), .G(I_1039_D), .S(I_2071_S));
  generic_nmos I_1136(.D(I_1136_D), .G(I_1137_G), .S(I_1168_D));
  generic_pmos I_1137(.D(I_1137_D), .G(I_1137_G), .S(I_1169_D));
  generic_nmos I_1138(.D(I_1139_D), .G(I_1269_S), .S(VSS));
  generic_pmos I_1139(.D(I_1139_D), .G(I_1269_S), .S(VDD));
  generic_nmos I_114(.D(I_114_D), .G(I_114_G), .S(I_146_D));
  generic_nmos I_1140(.D(I_1237_D), .G(I_1205_D), .S(VSS));
  generic_pmos I_1141(.D(I_1237_D), .G(I_1205_D), .S(VDD));
  generic_nmos I_1142(.D(I_1239_D), .G(I_1207_D), .S(VSS));
  generic_pmos I_1143(.D(I_1239_D), .G(I_1207_D), .S(VDD));
  generic_nmos I_1144(.D(I_1144_D), .G(I_1145_G), .S(VSS));
  generic_pmos I_1145(.D(I_1145_D), .G(I_1145_G), .S(VDD));
  generic_nmos I_1146(.D(I_1211_D), .G(I_735_D), .S(I_1178_D));
  generic_pmos I_1147(.D(I_1211_D), .G(I_735_D), .S(VDD));
  generic_nmos I_1148(.D(I_1213_D), .G(I_957_S), .S(I_1180_D));
  generic_pmos I_1149(.D(I_1213_D), .G(I_957_S), .S(VDD));
  generic_pmos I_115(.D(I_115_D), .G(I_146_G), .S(I_147_D));
  generic_nmos I_1150(.D(I_1279_S), .G(I_1119_D), .S(VSS));
  generic_pmos I_1151(.D(I_1279_S), .G(I_1119_D), .S(VDD));
  generic_nmos I_1152(.D(VSS), .G(I_1153_G), .S(I_1184_D));
  generic_pmos I_1153(.D(VDD), .G(I_1153_G), .S(I_1185_D));
  generic_nmos I_1154(.D(I_1187_S), .G(I_1539_D), .S(VSS));
  generic_pmos I_1155(.D(I_1187_S), .G(I_1539_D), .S(VDD));
  generic_nmos I_1156(.D(VSS), .G(I_1187_S), .S(I_1188_D));
  generic_pmos I_1157(.D(VDD), .G(I_1187_S), .S(I_1189_D));
  generic_nmos I_1158(.D(I_1158_D), .G(I_1253_S), .S(VSS));
  generic_pmos I_1159(.D(I_1223_D), .G(I_1253_S), .S(VDD));
  generic_nmos I_116(.D(I_116_D), .G(I_116_G), .S(I_148_D));
  generic_nmos I_1160(.D(VSS), .G(I_1193_G), .S(I_1259_S));
  generic_pmos I_1161(.D(VDD), .G(I_1193_G), .S(I_1259_S));
  generic_nmos I_1162(.D(VSS), .G(I_1259_D), .S(I_1195_D));
  generic_pmos I_1163(.D(VDD), .G(I_1259_D), .S(I_1195_D));
  generic_nmos I_1164(.D(I_1164_D), .G(I_1165_G), .S(I_1196_D));
  generic_pmos I_1165(.D(I_1165_D), .G(I_1165_G), .S(I_1197_D));
  generic_nmos I_1166(.D(I_1166_D), .G(I_1103_D), .S(I_2071_S));
  generic_pmos I_1167(.D(I_2071_S), .G(I_1103_D), .S(VDD));
  generic_nmos I_1168(.D(I_1168_D), .G(I_1169_G), .S(I_1200_D));
  generic_pmos I_1169(.D(I_1169_D), .G(I_1169_G), .S(I_1201_D));
  generic_pmos I_117(.D(I_117_D), .G(I_148_G), .S(I_149_D));
  generic_nmos I_1170(.D(VSS), .G(I_1267_D), .S(I_1269_S));
  generic_pmos I_1171(.D(VDD), .G(I_1267_D), .S(I_1269_S));
  generic_nmos I_1172(.D(VSS), .G(I_1269_D), .S(I_1205_D));
  generic_pmos I_1173(.D(VDD), .G(I_1269_D), .S(I_1205_D));
  generic_nmos I_1174(.D(VSS), .G(I_1271_D), .S(I_1207_D));
  generic_pmos I_1175(.D(VDD), .G(I_1271_D), .S(I_1207_D));
  generic_nmos I_1176(.D(VSS), .G(I_1435_D), .S(I_1208_D));
  generic_pmos I_1177(.D(VDD), .G(I_1435_D), .S(I_1209_D));
  generic_nmos I_1178(.D(I_1178_D), .G(I_1051_S), .S(I_1210_D));
  generic_pmos I_1179(.D(VDD), .G(I_1051_S), .S(I_1211_D));
  generic_nmos I_118(.D(I_118_D), .G(I_118_G), .S(I_151_D));
  generic_nmos I_1180(.D(I_1180_D), .G(I_511_D), .S(I_1212_D));
  generic_pmos I_1181(.D(VDD), .G(I_511_D), .S(I_1213_D));
  generic_nmos I_1182(.D(VSS), .G(I_1183_G), .S(VSS));
  generic_pmos I_1183(.D(VDD), .G(I_1183_G), .S(VDD));
  generic_nmos I_1184(.D(I_1184_D), .G(I_1185_G), .S(I_1185_D));
  generic_pmos I_1185(.D(I_1185_D), .G(I_1185_G), .S(VDD));
  generic_nmos I_1186(.D(VSS), .G(I_1539_D), .S(I_1187_S));
  generic_pmos I_1187(.D(VDD), .G(I_1539_D), .S(I_1187_S));
  generic_nmos I_1188(.D(I_1188_D), .G(I_1253_D), .S(I_1189_D));
  generic_pmos I_1189(.D(I_1189_D), .G(I_1253_D), .S(VDD));
  generic_pmos I_119(.D(VDD), .G(I_151_G), .S(I_151_D));
  generic_nmos I_1190(.D(VSS), .G(I_1255_D), .S(I_1253_S));
  generic_pmos I_1191(.D(VDD), .G(I_1255_D), .S(I_1253_S));
  generic_nmos I_1192(.D(I_1259_S), .G(I_1193_G), .S(VSS));
  generic_pmos I_1193(.D(I_1259_S), .G(I_1193_G), .S(VDD));
  generic_nmos I_1194(.D(I_1195_D), .G(I_1259_D), .S(VSS));
  generic_pmos I_1195(.D(I_1195_D), .G(I_1259_D), .S(VDD));
  generic_nmos I_1196(.D(I_1196_D), .G(I_1197_G), .S(I_1196_S));
  generic_pmos I_1197(.D(I_1197_D), .G(I_1197_G), .S(I_1197_S));
  generic_nmos I_1198(.D(I_2071_S), .G(I_1199_G), .S(I_1198_S));
  generic_pmos I_1199(.D(VDD), .G(I_1199_G), .S(I_1199_S));
  generic_nmos I_12(.D(I_12_D), .G(I_13_G), .S(I_44_D));
  generic_nmos I_120(.D(I_155_D), .G(I_315_D), .S(I_153_D));
  generic_nmos I_1200(.D(I_1200_D), .G(I_1201_G), .S(I_1200_S));
  generic_pmos I_1201(.D(I_1201_D), .G(I_1201_G), .S(I_1201_S));
  generic_nmos I_1202(.D(I_1269_S), .G(I_1267_D), .S(VSS));
  generic_pmos I_1203(.D(I_1269_S), .G(I_1267_D), .S(VDD));
  generic_nmos I_1204(.D(I_1205_D), .G(I_1269_D), .S(VSS));
  generic_pmos I_1205(.D(I_1205_D), .G(I_1269_D), .S(VDD));
  generic_nmos I_1206(.D(I_1207_D), .G(I_1271_D), .S(VSS));
  generic_pmos I_1207(.D(I_1207_D), .G(I_1271_D), .S(VDD));
  generic_nmos I_1208(.D(I_1208_D), .G(I_1435_D), .S(I_1209_S));
  generic_pmos I_1209(.D(I_1209_D), .G(I_1435_D), .S(I_1209_S));
  generic_pmos I_121(.D(I_155_D), .G(I_251_S), .S(I_153_D));
  generic_nmos I_1210(.D(I_1210_D), .G(I_1397_D), .S(VSS));
  generic_pmos I_1211(.D(I_1211_D), .G(I_1397_D), .S(VDD));
  generic_nmos I_1212(.D(I_1212_D), .G(I_477_S), .S(VSS));
  generic_pmos I_1213(.D(I_1213_D), .G(I_477_S), .S(VDD));
  generic_nmos I_1214(.D(VSS), .G(I_1279_S), .S(I_1247_D));
  generic_pmos I_1215(.D(VDD), .G(I_1279_S), .S(I_1247_D));
  generic_nmos I_1216(.D(VSS), .G(I_1251_D), .S(I_1249_D));
  generic_pmos I_1217(.D(VDD), .G(I_1251_D), .S(I_1249_D));
  generic_nmos I_1218(.D(I_1251_D), .G(I_1091_D), .S(I_1250_D));
  generic_pmos I_1219(.D(VDD), .G(I_1250_G), .S(I_1251_D));
  generic_nmos I_122(.D(I_2041_D), .G(I_1045_D), .S(I_155_D));
  generic_nmos I_1220(.D(I_1221_D), .G(I_1097_S), .S(I_1253_D));
  generic_pmos I_1221(.D(I_1221_D), .G(I_715_D), .S(I_1253_D));
  generic_nmos I_1222(.D(I_1223_D), .G(I_715_D), .S(I_1255_D));
  generic_pmos I_1223(.D(I_1223_D), .G(I_1097_S), .S(I_1255_D));
  generic_nmos I_1224(.D(I_1225_D), .G(I_1258_G), .S(I_1257_D));
  generic_pmos I_1225(.D(I_1225_D), .G(I_1099_S), .S(I_1257_D));
  generic_nmos I_1226(.D(I_1227_D), .G(I_1099_S), .S(I_1259_D));
  generic_pmos I_1227(.D(I_1227_D), .G(I_1258_G), .S(I_1259_D));
  generic_nmos I_1228(.D(I_1228_D), .G(I_1228_G), .S(VSS));
  generic_pmos I_1229(.D(I_1417_S), .G(I_1260_G), .S(VDD));
  generic_pmos I_123(.D(I_2041_D), .G(I_789_D), .S(I_155_D));
  generic_nmos I_1230(.D(I_1230_D), .G(I_1230_G), .S(VSS));
  generic_pmos I_1231(.D(I_1267_S), .G(I_1262_G), .S(VDD));
  generic_nmos I_1232(.D(I_1361_S), .G(I_1999_D), .S(I_1265_D));
  generic_pmos I_1233(.D(I_1361_S), .G(I_1297_D), .S(I_1265_D));
  generic_nmos I_1234(.D(I_1235_D), .G(I_735_D), .S(I_1267_D));
  generic_pmos I_1235(.D(I_1235_D), .G(I_1301_D), .S(I_1267_D));
  generic_nmos I_1236(.D(I_1237_D), .G(I_1301_D), .S(I_1269_D));
  generic_pmos I_1237(.D(I_1237_D), .G(I_735_D), .S(I_1269_D));
  generic_nmos I_1238(.D(I_1239_D), .G(I_315_D), .S(I_1271_D));
  generic_pmos I_1239(.D(I_1239_D), .G(I_251_S), .S(I_1271_D));
  generic_nmos I_124(.D(I_477_D), .G(I_93_S), .S(I_157_D));
  generic_nmos I_1240(.D(VSS), .G(I_1209_S), .S(I_1272_D));
  generic_pmos I_1241(.D(VDD), .G(I_1209_S), .S(I_1273_D));
  generic_nmos I_1242(.D(I_1275_D), .G(I_1307_D), .S(I_1274_D));
  generic_pmos I_1243(.D(VDD), .G(I_735_D), .S(I_1275_D));
  generic_nmos I_1244(.D(I_1244_D), .G(I_1244_G), .S(VSS));
  generic_pmos I_1245(.D(I_1407_D), .G(I_1343_D), .S(VDD));
  generic_nmos I_1246(.D(I_1247_D), .G(I_1469_D), .S(I_1279_D));
  generic_pmos I_1247(.D(I_1247_D), .G(I_1213_D), .S(I_1279_D));
  generic_nmos I_1248(.D(I_1249_D), .G(I_1251_D), .S(VSS));
  generic_pmos I_1249(.D(I_1249_D), .G(I_1251_D), .S(VDD));
  generic_pmos I_125(.D(I_477_D), .G(I_95_D), .S(I_157_D));
  generic_nmos I_1250(.D(I_1250_D), .G(I_1250_G), .S(VSS));
  generic_pmos I_1251(.D(I_1251_D), .G(I_1091_D), .S(VDD));
  generic_nmos I_1252(.D(I_1253_D), .G(I_715_D), .S(I_1253_S));
  generic_pmos I_1253(.D(I_1253_D), .G(I_1097_S), .S(I_1253_S));
  generic_nmos I_1254(.D(I_1255_D), .G(I_1097_S), .S(I_2329_D));
  generic_pmos I_1255(.D(I_1255_D), .G(I_715_D), .S(I_2329_D));
  generic_nmos I_1256(.D(I_1257_D), .G(I_1099_S), .S(I_1355_D));
  generic_pmos I_1257(.D(I_1257_D), .G(I_1258_G), .S(I_1355_D));
  generic_nmos I_1258(.D(I_1259_D), .G(I_1258_G), .S(I_1259_S));
  generic_pmos I_1259(.D(I_1259_D), .G(I_1099_S), .S(I_1259_S));
  generic_nmos I_126(.D(I_1407_D), .G(I_93_S), .S(I_159_S));
  generic_nmos I_1260(.D(VSS), .G(I_1260_G), .S(I_1417_S));
  generic_pmos I_1261(.D(VDD), .G(I_1261_G), .S(I_1261_S));
  generic_nmos I_1262(.D(VSS), .G(I_1262_G), .S(I_1267_S));
  generic_pmos I_1263(.D(VDD), .G(I_1263_G), .S(I_1263_S));
  generic_nmos I_1264(.D(I_1265_D), .G(I_1297_D), .S(I_2071_S));
  generic_pmos I_1265(.D(I_1265_D), .G(I_1999_D), .S(I_2071_S));
  generic_nmos I_1266(.D(I_1267_D), .G(I_1301_D), .S(I_1267_S));
  generic_pmos I_1267(.D(I_1267_D), .G(I_735_D), .S(I_1267_S));
  generic_nmos I_1268(.D(I_1269_D), .G(I_735_D), .S(I_1269_S));
  generic_pmos I_1269(.D(I_1269_D), .G(I_1301_D), .S(I_1269_S));
  generic_pmos I_127(.D(I_127_D), .G(I_158_G), .S(I_1407_D));
  generic_nmos I_1270(.D(I_1271_D), .G(I_251_S), .S(I_1335_D));
  generic_pmos I_1271(.D(I_1271_D), .G(I_315_D), .S(I_1335_D));
  generic_nmos I_1272(.D(I_1272_D), .G(I_1209_S), .S(I_1273_S));
  generic_pmos I_1273(.D(I_1273_D), .G(I_1209_S), .S(I_1273_S));
  generic_nmos I_1274(.D(I_1274_D), .G(I_735_D), .S(VSS));
  generic_pmos I_1275(.D(I_1275_D), .G(I_1307_D), .S(VDD));
  generic_nmos I_1276(.D(VSS), .G(I_1343_D), .S(I_1407_D));
  generic_pmos I_1277(.D(VDD), .G(I_1343_D), .S(I_1407_D));
  generic_nmos I_1278(.D(I_1279_D), .G(I_1213_D), .S(I_1279_S));
  generic_pmos I_1279(.D(I_1279_D), .G(I_1469_D), .S(I_1279_S));
  generic_nmos I_128(.D(I_128_D), .G(I_1089_D), .S(VSS));
  generic_nmos I_1280(.D(I_1280_D), .G(I_1281_G), .S(VSS));
  generic_pmos I_1281(.D(I_1281_D), .G(I_1281_G), .S(VDD));
  generic_nmos I_1282(.D(I_1283_D), .G(I_1345_D), .S(VSS));
  generic_pmos I_1283(.D(I_1283_D), .G(I_1345_D), .S(VDD));
  generic_nmos I_1284(.D(I_1381_D), .G(I_1349_D), .S(VSS));
  generic_pmos I_1285(.D(I_1381_D), .G(I_1349_D), .S(VDD));
  generic_nmos I_1286(.D(I_1383_D), .G(I_1187_S), .S(I_1318_D));
  generic_pmos I_1287(.D(VDD), .G(I_1187_S), .S(I_1383_D));
  generic_nmos I_1288(.D(I_1385_D), .G(I_1419_S), .S(VSS));
  generic_pmos I_1289(.D(I_1385_D), .G(I_1419_S), .S(VDD));
  generic_pmos I_129(.D(I_129_D), .G(I_225_D), .S(VDD));
  generic_nmos I_1290(.D(I_1387_D), .G(I_1355_D), .S(VSS));
  generic_pmos I_1291(.D(I_1387_D), .G(I_1355_D), .S(VDD));
  generic_nmos I_1292(.D(I_1292_D), .G(I_1293_G), .S(I_1324_D));
  generic_pmos I_1293(.D(I_1293_D), .G(I_1293_G), .S(I_1325_D));
  generic_nmos I_1294(.D(I_1295_D), .G(I_1997_D), .S(VSS));
  generic_pmos I_1295(.D(I_1295_D), .G(I_1997_D), .S(VDD));
  generic_nmos I_1296(.D(I_1297_D), .G(I_1999_D), .S(VSS));
  generic_pmos I_1297(.D(I_1297_D), .G(I_1999_D), .S(VDD));
  generic_nmos I_1298(.D(I_1298_D), .G(I_1299_G), .S(I_1331_D));
  generic_pmos I_1299(.D(I_1299_D), .G(I_1299_G), .S(I_1331_D));
  generic_pmos I_13(.D(I_13_D), .G(I_13_G), .S(I_45_D));
  generic_nmos I_130(.D(VSS), .G(I_130_G), .S(I_130_S));
  generic_nmos I_1300(.D(I_1301_D), .G(I_735_D), .S(VSS));
  generic_pmos I_1301(.D(I_1301_D), .G(I_735_D), .S(VDD));
  generic_nmos I_1302(.D(VSS), .G(I_1431_D), .S(I_1335_D));
  generic_pmos I_1303(.D(VDD), .G(I_1431_D), .S(I_1335_D));
  generic_nmos I_1304(.D(I_1304_D), .G(I_1305_G), .S(VSS));
  generic_pmos I_1305(.D(I_1305_D), .G(I_1305_G), .S(VDD));
  generic_nmos I_1306(.D(I_1307_D), .G(I_957_S), .S(VSS));
  generic_pmos I_1307(.D(I_1307_D), .G(I_957_S), .S(VDD));
  generic_nmos I_1308(.D(I_1309_D), .G(I_1369_S), .S(I_1340_D));
  generic_pmos I_1309(.D(I_1309_D), .G(I_1369_S), .S(I_1341_D));
  generic_pmos I_131(.D(VDD), .G(I_67_S), .S(I_131_S));
  generic_nmos I_1310(.D(I_1343_D), .G(I_1311_G), .S(I_1342_D));
  generic_pmos I_1311(.D(VDD), .G(I_1311_G), .S(I_1343_D));
  generic_nmos I_1312(.D(VSS), .G(I_1313_G), .S(I_1344_D));
  generic_pmos I_1313(.D(VDD), .G(I_1313_G), .S(I_1345_D));
  generic_nmos I_1314(.D(VSS), .G(I_1345_D), .S(I_1347_D));
  generic_pmos I_1315(.D(VDD), .G(I_1345_D), .S(I_1347_D));
  generic_nmos I_1316(.D(VSS), .G(I_1187_S), .S(I_1348_D));
  generic_pmos I_1317(.D(VDD), .G(I_1187_S), .S(I_1349_D));
  generic_nmos I_1318(.D(I_1318_D), .G(I_1413_S), .S(VSS));
  generic_pmos I_1319(.D(I_1383_D), .G(I_1413_S), .S(VDD));
  generic_nmos I_132(.D(I_133_D), .G(I_395_D), .S(I_133_S));
  generic_nmos I_1320(.D(VSS), .G(I_1417_D), .S(I_1419_S));
  generic_pmos I_1321(.D(VDD), .G(I_1417_D), .S(I_1419_S));
  generic_nmos I_1322(.D(VSS), .G(I_1419_D), .S(I_1355_D));
  generic_pmos I_1323(.D(VDD), .G(I_1419_D), .S(I_1355_D));
  generic_nmos I_1324(.D(I_1324_D), .G(I_1325_G), .S(I_1356_D));
  generic_pmos I_1325(.D(I_1325_D), .G(I_1325_G), .S(I_1357_D));
  generic_nmos I_1326(.D(VSS), .G(I_1997_D), .S(I_1358_D));
  generic_pmos I_1327(.D(VDD), .G(I_1997_D), .S(I_1359_D));
  generic_nmos I_1328(.D(VSS), .G(I_1329_G), .S(VSS));
  generic_pmos I_1329(.D(VDD), .G(I_1329_G), .S(VDD));
  generic_pmos I_133(.D(I_133_D), .G(I_329_D), .S(I_133_S));
  generic_nmos I_1330(.D(I_1331_D), .G(I_1365_S), .S(I_1362_D));
  generic_pmos I_1331(.D(I_1331_D), .G(I_1365_S), .S(I_1363_D));
  generic_nmos I_1332(.D(VSS), .G(I_1523_S), .S(I_1364_D));
  generic_pmos I_1333(.D(VDD), .G(I_1523_S), .S(I_1365_D));
  generic_nmos I_1334(.D(I_1335_D), .G(I_1431_D), .S(VSS));
  generic_pmos I_1335(.D(I_1335_D), .G(I_1431_D), .S(VDD));
  generic_nmos I_1336(.D(VSS), .G(I_1273_S), .S(I_1368_D));
  generic_pmos I_1337(.D(VDD), .G(I_1273_S), .S(I_1369_D));
  generic_nmos I_1338(.D(VSS), .G(I_1307_D), .S(I_1435_D));
  generic_pmos I_1339(.D(VDD), .G(I_1307_D), .S(I_1371_D));
  generic_nmos I_134(.D(I_135_D), .G(I_329_D), .S(I_2169_D));
  generic_nmos I_1340(.D(I_1340_D), .G(I_1369_S), .S(VSS));
  generic_pmos I_1341(.D(I_1341_D), .G(I_1369_S), .S(VDD));
  generic_nmos I_1342(.D(I_1342_D), .G(I_1439_D), .S(VSS));
  generic_pmos I_1343(.D(I_1343_D), .G(I_1439_D), .S(VDD));
  generic_nmos I_1344(.D(I_1344_D), .G(I_1409_D), .S(I_1345_D));
  generic_pmos I_1345(.D(I_1345_D), .G(I_1409_D), .S(VDD));
  generic_nmos I_1346(.D(I_1347_D), .G(I_1345_D), .S(VSS));
  generic_pmos I_1347(.D(I_1347_D), .G(I_1345_D), .S(VDD));
  generic_nmos I_1348(.D(I_1348_D), .G(I_1413_D), .S(I_1349_D));
  generic_pmos I_1349(.D(I_1349_D), .G(I_1413_D), .S(VDD));
  generic_pmos I_135(.D(I_135_D), .G(I_395_D), .S(I_2169_D));
  generic_nmos I_1350(.D(VSS), .G(I_1415_D), .S(I_1413_S));
  generic_pmos I_1351(.D(VDD), .G(I_1415_D), .S(I_1413_S));
  generic_nmos I_1352(.D(I_1419_S), .G(I_1417_D), .S(VSS));
  generic_pmos I_1353(.D(I_1419_S), .G(I_1417_D), .S(VDD));
  generic_nmos I_1354(.D(I_1355_D), .G(I_1419_D), .S(VSS));
  generic_pmos I_1355(.D(I_1355_D), .G(I_1419_D), .S(VDD));
  generic_nmos I_1356(.D(I_1356_D), .G(I_1357_G), .S(I_1356_S));
  generic_pmos I_1357(.D(I_1357_D), .G(I_1357_G), .S(I_1357_S));
  generic_nmos I_1358(.D(I_1358_D), .G(I_3111_S), .S(I_1359_D));
  generic_pmos I_1359(.D(I_1359_D), .G(I_3111_S), .S(VDD));
  generic_nmos I_136(.D(I_136_D), .G(I_136_G), .S(I_136_S));
  generic_nmos I_1360(.D(VSS), .G(I_2071_S), .S(I_1361_S));
  generic_pmos I_1361(.D(VDD), .G(I_2071_S), .S(I_1361_S));
  generic_nmos I_1362(.D(I_1362_D), .G(I_1365_S), .S(VSS));
  generic_pmos I_1363(.D(I_1363_D), .G(I_1365_S), .S(VDD));
  generic_nmos I_1364(.D(I_1364_D), .G(I_1523_S), .S(I_1365_S));
  generic_pmos I_1365(.D(I_1365_D), .G(I_1523_S), .S(I_1365_S));
  generic_nmos I_1366(.D(VSS), .G(I_1335_D), .S(I_1399_D));
  generic_pmos I_1367(.D(VDD), .G(I_1335_D), .S(I_1399_D));
  generic_nmos I_1368(.D(I_1368_D), .G(I_1273_S), .S(I_1369_S));
  generic_pmos I_1369(.D(I_1369_D), .G(I_1273_S), .S(I_1369_S));
  generic_pmos I_137(.D(I_137_D), .G(I_137_G), .S(I_137_S));
  generic_nmos I_1370(.D(I_1435_D), .G(I_1051_S), .S(VSS));
  generic_pmos I_1371(.D(I_1371_D), .G(I_1051_S), .S(I_1403_D));
  generic_nmos I_1372(.D(VSS), .G(I_1247_D), .S(I_1373_S));
  generic_pmos I_1373(.D(VDD), .G(I_1247_D), .S(I_1373_S));
  generic_nmos I_1374(.D(VSS), .G(I_1375_G), .S(I_1374_S));
  generic_pmos I_1375(.D(VDD), .G(I_1375_G), .S(I_1375_S));
  generic_nmos I_1376(.D(I_1409_D), .G(I_1409_G), .S(I_1408_D));
  generic_pmos I_1377(.D(VDD), .G(I_1408_G), .S(I_1409_D));
  generic_nmos I_1378(.D(I_1411_S), .G(I_1671_S), .S(VSS));
  generic_pmos I_1379(.D(I_1379_D), .G(I_1410_G), .S(VDD));
  generic_nmos I_138(.D(I_138_D), .G(I_138_G), .S(I_138_S));
  generic_nmos I_1380(.D(I_1381_D), .G(I_1097_S), .S(I_1413_D));
  generic_pmos I_1381(.D(I_1381_D), .G(I_715_D), .S(I_1413_D));
  generic_nmos I_1382(.D(I_1383_D), .G(I_715_D), .S(I_1415_D));
  generic_pmos I_1383(.D(I_1383_D), .G(I_1097_S), .S(I_1415_D));
  generic_nmos I_1384(.D(I_1385_D), .G(I_1101_S), .S(I_1417_D));
  generic_pmos I_1385(.D(I_1385_D), .G(I_1420_S), .S(I_1417_D));
  generic_nmos I_1386(.D(I_1387_D), .G(I_1420_S), .S(I_1419_D));
  generic_pmos I_1387(.D(I_1387_D), .G(I_1101_S), .S(I_1419_D));
  generic_nmos I_1388(.D(I_1388_D), .G(I_1388_G), .S(VSS));
  generic_pmos I_1389(.D(I_1420_S), .G(I_1101_S), .S(VDD));
  generic_pmos I_139(.D(I_139_D), .G(I_139_G), .S(I_139_S));
  generic_nmos I_1390(.D(VSS), .G(I_1295_D), .S(I_1422_D));
  generic_pmos I_1391(.D(VDD), .G(I_2631_S), .S(I_1423_D));
  generic_nmos I_1392(.D(I_1999_D), .G(I_2071_S), .S(I_1425_S));
  generic_pmos I_1393(.D(I_1393_D), .G(I_1361_S), .S(I_1999_D));
  generic_nmos I_1394(.D(I_1525_D), .G(I_1589_S), .S(I_1427_D));
  generic_pmos I_1395(.D(I_1525_D), .G(I_1749_S), .S(I_1427_D));
  generic_nmos I_1396(.D(I_1397_D), .G(I_1749_S), .S(I_1429_D));
  generic_pmos I_1397(.D(I_1397_D), .G(I_1589_S), .S(I_1429_D));
  generic_nmos I_1398(.D(I_1399_D), .G(I_251_S), .S(I_1431_D));
  generic_pmos I_1399(.D(I_1399_D), .G(I_315_D), .S(I_1431_D));
  generic_nmos I_14(.D(I_14_D), .G(I_15_G), .S(I_46_D));
  generic_nmos I_140(.D(I_140_D), .G(I_140_G), .S(I_140_S));
  generic_nmos I_1400(.D(I_1401_D), .G(I_789_D), .S(I_1433_D));
  generic_pmos I_1401(.D(I_1401_D), .G(I_1045_D), .S(I_1433_D));
  generic_nmos I_1402(.D(I_1402_D), .G(I_1402_G), .S(VSS));
  generic_pmos I_1403(.D(I_1403_D), .G(I_1373_S), .S(I_1435_D));
  generic_nmos I_1404(.D(VSS), .G(I_1397_D), .S(I_1913_S));
  generic_pmos I_1405(.D(VDD), .G(I_735_D), .S(I_1437_D));
  generic_nmos I_1406(.D(I_1407_D), .G(I_93_S), .S(I_1439_D));
  generic_pmos I_1407(.D(I_1407_D), .G(I_95_D), .S(I_1439_D));
  generic_nmos I_1408(.D(I_1408_D), .G(I_1408_G), .S(VSS));
  generic_pmos I_1409(.D(I_1409_D), .G(I_1409_G), .S(VDD));
  generic_pmos I_141(.D(I_141_D), .G(I_141_G), .S(I_141_S));
  generic_nmos I_1410(.D(VSS), .G(I_1410_G), .S(I_1410_S));
  generic_pmos I_1411(.D(VDD), .G(I_1671_S), .S(I_1411_S));
  generic_nmos I_1412(.D(I_1413_D), .G(I_715_D), .S(I_1413_S));
  generic_pmos I_1413(.D(I_1413_D), .G(I_1097_S), .S(I_1413_S));
  generic_nmos I_1414(.D(I_1415_D), .G(I_1097_S), .S(I_1415_S));
  generic_pmos I_1415(.D(I_1415_D), .G(I_715_D), .S(I_1415_S));
  generic_nmos I_1416(.D(I_1417_D), .G(I_1420_S), .S(I_1417_S));
  generic_pmos I_1417(.D(I_1417_D), .G(I_1101_S), .S(I_1417_S));
  generic_nmos I_1418(.D(I_1419_D), .G(I_1101_S), .S(I_1419_S));
  generic_pmos I_1419(.D(I_1419_D), .G(I_1420_S), .S(I_1419_S));
  generic_nmos I_142(.D(I_142_D), .G(I_142_G), .S(I_142_S));
  generic_nmos I_1420(.D(VSS), .G(I_1101_S), .S(I_1420_S));
  generic_pmos I_1421(.D(VDD), .G(I_1421_G), .S(I_1421_S));
  generic_nmos I_1422(.D(I_1422_D), .G(I_2631_S), .S(I_1423_D));
  generic_pmos I_1423(.D(I_1423_D), .G(I_1295_D), .S(VDD));
  generic_nmos I_1424(.D(I_1425_S), .G(I_1361_S), .S(VSS));
  generic_pmos I_1425(.D(I_1999_D), .G(I_1361_S), .S(I_1425_S));
  generic_nmos I_1426(.D(I_1427_D), .G(I_1749_S), .S(I_1523_S));
  generic_pmos I_1427(.D(I_1427_D), .G(I_1589_S), .S(I_1523_S));
  generic_nmos I_1428(.D(I_1429_D), .G(I_1589_S), .S(I_1461_D));
  generic_pmos I_1429(.D(I_1429_D), .G(I_1749_S), .S(I_1461_D));
  generic_pmos I_143(.D(I_143_D), .G(I_143_G), .S(I_143_S));
  generic_nmos I_1430(.D(I_1431_D), .G(I_315_D), .S(I_1433_D));
  generic_pmos I_1431(.D(I_1431_D), .G(I_251_S), .S(I_1433_D));
  generic_nmos I_1432(.D(I_1433_D), .G(I_1045_D), .S(I_2521_D));
  generic_pmos I_1433(.D(I_1433_D), .G(I_789_D), .S(I_2521_D));
  generic_nmos I_1434(.D(VSS), .G(I_1373_S), .S(I_1435_D));
  generic_pmos I_1435(.D(I_1435_D), .G(I_1435_G), .S(I_1435_S));
  generic_nmos I_1436(.D(I_1913_S), .G(I_735_D), .S(VSS));
  generic_pmos I_1437(.D(I_1437_D), .G(I_1397_D), .S(I_1913_S));
  generic_nmos I_1438(.D(I_1439_D), .G(I_95_D), .S(I_1439_S));
  generic_pmos I_1439(.D(I_1439_D), .G(I_93_S), .S(I_1439_S));
  generic_nmos I_144(.D(I_144_D), .G(I_144_G), .S(I_144_S));
  generic_nmos I_1440(.D(I_1537_D), .G(I_1571_S), .S(VSS));
  generic_pmos I_1441(.D(I_1537_D), .G(I_1571_S), .S(VDD));
  generic_nmos I_1442(.D(I_1539_D), .G(I_1507_D), .S(VSS));
  generic_pmos I_1443(.D(I_1539_D), .G(I_1507_D), .S(VDD));
  generic_nmos I_1444(.D(I_1541_D), .G(I_1575_S), .S(VSS));
  generic_pmos I_1445(.D(I_1541_D), .G(I_1575_S), .S(VDD));
  generic_nmos I_1446(.D(I_1573_S), .G(I_1511_S), .S(I_1478_D));
  generic_pmos I_1447(.D(VDD), .G(I_1511_S), .S(I_1573_S));
  generic_nmos I_1448(.D(I_1448_D), .G(I_1449_G), .S(I_1480_D));
  generic_pmos I_1449(.D(I_1449_D), .G(I_1449_G), .S(I_1481_D));
  generic_pmos I_145(.D(I_145_D), .G(I_145_G), .S(I_145_S));
  generic_nmos I_1450(.D(I_1483_D), .G(I_1195_D), .S(I_1482_D));
  generic_pmos I_1451(.D(VDD), .G(I_1195_D), .S(I_1483_D));
  generic_nmos I_1452(.D(I_1452_D), .G(I_1453_G), .S(I_1484_D));
  generic_pmos I_1453(.D(I_1453_D), .G(I_1453_G), .S(I_1485_D));
  generic_nmos I_1454(.D(VSS), .G(I_1359_D), .S(I_1486_D));
  generic_pmos I_1455(.D(VDD), .G(I_1359_D), .S(I_1518_D));
  generic_nmos I_1456(.D(I_1456_D), .G(I_1457_G), .S(I_1488_D));
  generic_pmos I_1457(.D(I_1457_D), .G(I_1457_G), .S(I_1489_D));
  generic_nmos I_1458(.D(VSS), .G(I_1427_D), .S(I_1491_D));
  generic_pmos I_1459(.D(VDD), .G(I_1427_D), .S(I_1491_D));
  generic_nmos I_146(.D(I_146_D), .G(I_146_G), .S(I_146_S));
  generic_nmos I_1460(.D(I_1461_D), .G(I_1525_D), .S(VSS));
  generic_pmos I_1461(.D(I_1461_D), .G(I_1525_D), .S(VDD));
  generic_nmos I_1462(.D(I_1559_D), .G(I_1593_S), .S(VSS));
  generic_pmos I_1463(.D(I_1559_D), .G(I_1593_S), .S(VDD));
  generic_nmos I_1464(.D(I_1561_D), .G(I_1529_D), .S(VSS));
  generic_pmos I_1465(.D(I_1561_D), .G(I_1529_D), .S(VDD));
  generic_nmos I_1466(.D(I_1499_D), .G(I_1051_S), .S(I_1498_D));
  generic_pmos I_1467(.D(VDD), .G(I_1051_S), .S(I_1499_D));
  generic_nmos I_1468(.D(I_1469_D), .G(I_1213_D), .S(VSS));
  generic_pmos I_1469(.D(I_1469_D), .G(I_1213_D), .S(VDD));
  generic_pmos I_147(.D(I_147_D), .G(I_147_G), .S(I_147_S));
  generic_nmos I_1470(.D(I_1535_D), .G(I_3667_D), .S(I_1502_D));
  generic_pmos I_1471(.D(I_1535_D), .G(I_3667_D), .S(VDD));
  generic_nmos I_1472(.D(VSS), .G(I_1569_D), .S(I_1571_S));
  generic_pmos I_1473(.D(VDD), .G(I_1569_D), .S(I_1571_S));
  generic_nmos I_1474(.D(VSS), .G(I_1571_D), .S(I_1507_D));
  generic_pmos I_1475(.D(VDD), .G(I_1571_D), .S(I_1507_D));
  generic_nmos I_1476(.D(VSS), .G(I_1347_D), .S(I_1508_D));
  generic_pmos I_1477(.D(VDD), .G(I_1347_D), .S(I_1575_S));
  generic_nmos I_1478(.D(I_1478_D), .G(I_1347_D), .S(VSS));
  generic_pmos I_1479(.D(I_1573_S), .G(I_1347_D), .S(VDD));
  generic_nmos I_148(.D(I_148_D), .G(I_148_G), .S(I_148_S));
  generic_nmos I_1480(.D(I_1480_D), .G(I_1481_G), .S(I_1512_D));
  generic_pmos I_1481(.D(I_1481_D), .G(I_1481_G), .S(I_1513_D));
  generic_nmos I_1482(.D(I_1482_D), .G(VDD), .S(VSS));
  generic_pmos I_1483(.D(I_1483_D), .G(VDD), .S(VDD));
  generic_nmos I_1484(.D(I_1484_D), .G(I_1485_G), .S(I_1516_D));
  generic_pmos I_1485(.D(I_1485_D), .G(I_1485_G), .S(I_1517_D));
  generic_nmos I_1486(.D(I_1486_D), .G(I_1423_D), .S(I_1518_D));
  generic_pmos I_1487(.D(I_1518_D), .G(I_1423_D), .S(VDD));
  generic_nmos I_1488(.D(I_1488_D), .G(I_1489_G), .S(I_1520_D));
  generic_pmos I_1489(.D(I_1489_D), .G(I_1489_G), .S(I_1521_D));
  generic_pmos I_149(.D(I_149_D), .G(I_149_G), .S(I_149_S));
  generic_nmos I_1490(.D(I_1491_D), .G(I_1427_D), .S(VSS));
  generic_pmos I_1491(.D(I_1491_D), .G(I_1427_D), .S(VDD));
  generic_nmos I_1492(.D(VSS), .G(I_1429_D), .S(I_1525_D));
  generic_pmos I_1493(.D(VDD), .G(I_1429_D), .S(I_1525_D));
  generic_nmos I_1494(.D(VSS), .G(I_1591_D), .S(I_1593_S));
  generic_pmos I_1495(.D(VDD), .G(I_1591_D), .S(I_1593_S));
  generic_nmos I_1496(.D(VSS), .G(I_1593_D), .S(I_1529_D));
  generic_pmos I_1497(.D(VDD), .G(I_1593_D), .S(I_1529_D));
  generic_nmos I_1498(.D(I_1498_D), .G(I_1997_D), .S(VSS));
  generic_pmos I_1499(.D(I_1499_D), .G(I_1997_D), .S(VDD));
  generic_pmos I_15(.D(I_15_D), .G(I_15_G), .S(I_47_D));
  generic_nmos I_150(.D(I_151_D), .G(I_151_G), .S(VSS));
  generic_nmos I_1500(.D(VSS), .G(I_1627_D), .S(I_1597_D));
  generic_pmos I_1501(.D(VDD), .G(I_1627_D), .S(I_1597_D));
  generic_nmos I_1502(.D(I_1502_D), .G(I_1758_S), .S(I_1534_D));
  generic_pmos I_1503(.D(VDD), .G(I_1758_S), .S(I_1535_D));
  generic_nmos I_1504(.D(I_1571_S), .G(I_1569_D), .S(VSS));
  generic_pmos I_1505(.D(I_1571_S), .G(I_1569_D), .S(VDD));
  generic_nmos I_1506(.D(I_1507_D), .G(I_1571_D), .S(VSS));
  generic_pmos I_1507(.D(I_1507_D), .G(I_1571_D), .S(VDD));
  generic_nmos I_1508(.D(I_1508_D), .G(I_1573_D), .S(I_1575_S));
  generic_pmos I_1509(.D(I_1575_S), .G(I_1573_D), .S(VDD));
  generic_pmos I_151(.D(I_151_D), .G(I_151_G), .S(VDD));
  generic_nmos I_1510(.D(VSS), .G(I_1575_D), .S(I_1511_S));
  generic_pmos I_1511(.D(VDD), .G(I_1575_D), .S(I_1511_S));
  generic_nmos I_1512(.D(I_1512_D), .G(I_1513_G), .S(I_1512_S));
  generic_pmos I_1513(.D(I_1513_D), .G(I_1513_G), .S(I_1513_S));
  generic_nmos I_1514(.D(VSS), .G(I_1483_D), .S(I_1515_S));
  generic_pmos I_1515(.D(VDD), .G(I_1483_D), .S(I_1515_S));
  generic_nmos I_1516(.D(I_1516_D), .G(I_1517_G), .S(I_1516_S));
  generic_pmos I_1517(.D(I_1517_D), .G(I_1517_G), .S(I_1517_S));
  generic_nmos I_1518(.D(I_1518_D), .G(I_1519_G), .S(I_1518_S));
  generic_pmos I_1519(.D(VDD), .G(I_1519_G), .S(I_1519_S));
  generic_nmos I_152(.D(I_153_D), .G(I_251_S), .S(I_185_D));
  generic_nmos I_1520(.D(I_1520_D), .G(I_1521_G), .S(I_1520_S));
  generic_pmos I_1521(.D(I_1521_D), .G(I_1521_G), .S(I_1521_S));
  generic_nmos I_1522(.D(VSS), .G(I_1491_D), .S(I_1523_S));
  generic_pmos I_1523(.D(VDD), .G(I_1491_D), .S(I_1523_S));
  generic_nmos I_1524(.D(I_1525_D), .G(I_1429_D), .S(VSS));
  generic_pmos I_1525(.D(I_1525_D), .G(I_1429_D), .S(VDD));
  generic_nmos I_1526(.D(I_1593_S), .G(I_1591_D), .S(VSS));
  generic_pmos I_1527(.D(I_1593_S), .G(I_1591_D), .S(VDD));
  generic_nmos I_1528(.D(I_1529_D), .G(I_1593_D), .S(VSS));
  generic_pmos I_1529(.D(I_1529_D), .G(I_1593_D), .S(VDD));
  generic_pmos I_153(.D(I_153_D), .G(I_315_D), .S(I_185_D));
  generic_nmos I_1530(.D(VSS), .G(I_1499_D), .S(I_1531_S));
  generic_pmos I_1531(.D(VDD), .G(I_1499_D), .S(I_1531_S));
  generic_nmos I_1532(.D(I_1597_D), .G(I_1627_D), .S(VSS));
  generic_pmos I_1533(.D(I_1597_D), .G(I_1627_D), .S(VDD));
  generic_nmos I_1534(.D(I_1534_D), .G(I_1598_S), .S(VSS));
  generic_pmos I_1535(.D(I_1535_D), .G(I_1598_S), .S(VDD));
  generic_nmos I_1536(.D(I_1537_D), .G(I_1671_S), .S(I_1569_D));
  generic_pmos I_1537(.D(I_1537_D), .G(I_1411_S), .S(I_1569_D));
  generic_nmos I_1538(.D(I_1539_D), .G(I_1411_S), .S(I_1571_D));
  generic_pmos I_1539(.D(I_1539_D), .G(I_1671_S), .S(I_1571_D));
  generic_nmos I_154(.D(I_155_D), .G(I_789_D), .S(VSS));
  generic_nmos I_1540(.D(I_1541_D), .G(I_1576_S), .S(I_1573_D));
  generic_pmos I_1541(.D(I_1541_D), .G(I_1051_S), .S(I_1573_D));
  generic_nmos I_1542(.D(I_1573_S), .G(I_1051_S), .S(I_1575_D));
  generic_pmos I_1543(.D(I_1573_S), .G(I_1576_S), .S(I_1575_D));
  generic_nmos I_1544(.D(I_1544_D), .G(I_1544_G), .S(VSS));
  generic_pmos I_1545(.D(I_1576_S), .G(I_1051_S), .S(VDD));
  generic_nmos I_1546(.D(I_1546_D), .G(I_1546_G), .S(I_1578_D));
  generic_pmos I_1547(.D(I_1547_D), .G(I_1578_G), .S(I_1579_D));
  generic_nmos I_1548(.D(I_1548_D), .G(I_1548_G), .S(I_1580_D));
  generic_pmos I_1549(.D(I_1549_D), .G(I_1580_G), .S(I_1581_D));
  generic_pmos I_155(.D(I_155_D), .G(I_1045_D), .S(VSS));
  generic_nmos I_1550(.D(I_1550_D), .G(I_1550_G), .S(I_1582_D));
  generic_pmos I_1551(.D(I_1551_D), .G(I_1582_G), .S(I_1583_D));
  generic_nmos I_1552(.D(I_1585_D), .G(I_1518_D), .S(I_1584_D));
  generic_pmos I_1553(.D(VDD), .G(I_1679_D), .S(I_1585_D));
  generic_nmos I_1554(.D(I_1554_D), .G(I_1554_G), .S(I_1586_D));
  generic_pmos I_1555(.D(I_1555_D), .G(I_1586_G), .S(I_1587_D));
  generic_nmos I_1556(.D(I_1589_S), .G(I_1588_S), .S(VSS));
  generic_pmos I_1557(.D(I_1588_S), .G(I_1685_D), .S(VDD));
  generic_nmos I_1558(.D(I_1559_D), .G(I_1623_D), .S(I_1591_D));
  generic_pmos I_1559(.D(I_1559_D), .G(I_1753_S), .S(I_1591_D));
  generic_nmos I_156(.D(I_157_D), .G(I_95_D), .S(I_253_S));
  generic_nmos I_1560(.D(I_1561_D), .G(I_1753_S), .S(I_1593_D));
  generic_pmos I_1561(.D(I_1561_D), .G(I_1623_D), .S(I_1593_D));
  generic_nmos I_1562(.D(VSS), .G(I_1531_S), .S(I_1627_D));
  generic_pmos I_1563(.D(VDD), .G(I_1531_S), .S(I_1627_D));
  generic_nmos I_1564(.D(VSS), .G(I_1627_D), .S(I_1597_D));
  generic_pmos I_1565(.D(VDD), .G(I_1627_D), .S(I_1597_D));
  generic_nmos I_1566(.D(I_1599_S), .G(I_1598_S), .S(VSS));
  generic_pmos I_1567(.D(I_1598_S), .G(I_1597_D), .S(VDD));
  generic_nmos I_1568(.D(I_1569_D), .G(I_1411_S), .S(I_1891_S));
  generic_pmos I_1569(.D(I_1569_D), .G(I_1671_S), .S(I_1891_S));
  generic_pmos I_157(.D(I_157_D), .G(I_93_S), .S(I_253_S));
  generic_nmos I_1570(.D(I_1571_D), .G(I_1671_S), .S(I_1571_S));
  generic_pmos I_1571(.D(I_1571_D), .G(I_1411_S), .S(I_1571_S));
  generic_nmos I_1572(.D(I_1573_D), .G(I_1051_S), .S(I_1573_S));
  generic_pmos I_1573(.D(I_1573_D), .G(I_1576_S), .S(I_1573_S));
  generic_nmos I_1574(.D(I_1575_D), .G(I_1576_S), .S(I_1575_S));
  generic_pmos I_1575(.D(I_1575_D), .G(I_1051_S), .S(I_1575_S));
  generic_nmos I_1576(.D(VSS), .G(I_1051_S), .S(I_1576_S));
  generic_pmos I_1577(.D(VDD), .G(I_1577_G), .S(I_1577_S));
  generic_nmos I_1578(.D(I_1578_D), .G(I_1578_G), .S(I_1578_S));
  generic_pmos I_1579(.D(I_1579_D), .G(I_1579_G), .S(I_1579_S));
  generic_nmos I_158(.D(I_159_S), .G(I_158_G), .S(I_158_S));
  generic_nmos I_1580(.D(I_1580_D), .G(I_1580_G), .S(I_1580_S));
  generic_pmos I_1581(.D(I_1581_D), .G(I_1581_G), .S(I_1581_S));
  generic_nmos I_1582(.D(I_1582_D), .G(I_1582_G), .S(I_1582_S));
  generic_pmos I_1583(.D(I_1583_D), .G(I_1583_G), .S(I_1583_S));
  generic_nmos I_1584(.D(I_1584_D), .G(I_1679_D), .S(VSS));
  generic_pmos I_1585(.D(I_1585_D), .G(I_1518_D), .S(VDD));
  generic_nmos I_1586(.D(I_1586_D), .G(I_1586_G), .S(I_1586_S));
  generic_pmos I_1587(.D(I_1587_D), .G(I_1587_G), .S(I_1587_S));
  generic_nmos I_1588(.D(VSS), .G(I_1685_D), .S(I_1588_S));
  generic_pmos I_1589(.D(VDD), .G(I_1588_S), .S(I_1589_S));
  generic_pmos I_159(.D(I_1407_D), .G(I_95_D), .S(I_159_S));
  generic_nmos I_1590(.D(I_1591_D), .G(I_1753_S), .S(I_1845_D));
  generic_pmos I_1591(.D(I_1591_D), .G(I_1623_D), .S(I_1845_D));
  generic_nmos I_1592(.D(I_1593_D), .G(I_1623_D), .S(I_1593_S));
  generic_pmos I_1593(.D(I_1593_D), .G(I_1753_S), .S(I_1593_S));
  generic_nmos I_1594(.D(I_1627_D), .G(I_1531_S), .S(VSS));
  generic_pmos I_1595(.D(I_1627_D), .G(I_1531_S), .S(VDD));
  generic_nmos I_1596(.D(I_1597_D), .G(I_1627_D), .S(VSS));
  generic_pmos I_1597(.D(I_1597_D), .G(I_1627_D), .S(VDD));
  generic_nmos I_1598(.D(VSS), .G(I_1597_D), .S(I_1598_S));
  generic_pmos I_1599(.D(VDD), .G(I_1598_S), .S(I_1599_S));
  generic_nmos I_16(.D(I_16_D), .G(I_17_G), .S(I_48_D));
  generic_nmos I_160(.D(I_224_D), .G(I_1832_D), .S(I_225_D));
  generic_nmos I_1600(.D(I_1697_D), .G(I_1731_S), .S(VSS));
  generic_pmos I_1601(.D(I_1697_D), .G(I_1731_S), .S(VDD));
  generic_nmos I_1602(.D(I_1699_D), .G(I_1667_D), .S(VSS));
  generic_pmos I_1603(.D(I_1699_D), .G(I_1667_D), .S(VDD));
  generic_nmos I_1604(.D(I_1701_D), .G(I_1735_S), .S(VSS));
  generic_pmos I_1605(.D(I_1701_D), .G(I_1735_S), .S(VDD));
  generic_nmos I_1606(.D(I_1733_S), .G(I_1671_S), .S(I_1638_D));
  generic_pmos I_1607(.D(VDD), .G(I_1671_S), .S(I_1733_S));
  generic_nmos I_1608(.D(I_1609_D), .G(I_1249_D), .S(VSS));
  generic_pmos I_1609(.D(I_1609_D), .G(I_1249_D), .S(VDD));
  generic_pmos I_161(.D(VDD), .G(I_1832_D), .S(I_193_D));
  generic_nmos I_1610(.D(I_1610_D), .G(I_1611_G), .S(I_1642_D));
  generic_pmos I_1611(.D(I_1611_D), .G(I_1611_G), .S(I_1643_D));
  generic_nmos I_1612(.D(I_1612_D), .G(I_1613_G), .S(I_1644_D));
  generic_pmos I_1613(.D(I_1613_D), .G(I_1613_G), .S(I_1645_D));
  generic_nmos I_1614(.D(I_1614_D), .G(I_1615_G), .S(VSS));
  generic_pmos I_1615(.D(I_1615_D), .G(I_1615_G), .S(VDD));
  generic_nmos I_1616(.D(VSS), .G(I_1518_D), .S(I_1648_D));
  generic_pmos I_1617(.D(I_1648_D), .G(I_1518_D), .S(I_1649_D));
  generic_nmos I_1618(.D(I_1618_D), .G(I_1619_G), .S(I_1650_D));
  generic_pmos I_1619(.D(I_1619_D), .G(I_1619_G), .S(I_1651_D));
  generic_nmos I_162(.D(I_162_D), .G(I_163_G), .S(VSS));
  generic_nmos I_1620(.D(I_1620_D), .G(I_1621_G), .S(VSS));
  generic_pmos I_1621(.D(I_1621_D), .G(I_1621_G), .S(VDD));
  generic_nmos I_1622(.D(I_1623_D), .G(I_1687_S), .S(VSS));
  generic_pmos I_1623(.D(I_1623_D), .G(I_1687_S), .S(VDD));
  generic_nmos I_1624(.D(I_1689_D), .G(I_1879_D), .S(VSS));
  generic_pmos I_1625(.D(I_1689_D), .G(I_1879_D), .S(VDD));
  generic_nmos I_1626(.D(I_1627_D), .G(I_1531_S), .S(VSS));
  generic_pmos I_1627(.D(I_1627_D), .G(I_1531_S), .S(VDD));
  generic_nmos I_1628(.D(I_1693_D), .G(I_1535_D), .S(I_1660_D));
  generic_pmos I_1629(.D(I_1693_D), .G(I_1535_D), .S(VDD));
  generic_pmos I_163(.D(I_163_D), .G(I_163_G), .S(VDD));
  generic_nmos I_1630(.D(I_1695_D), .G(I_1631_G), .S(I_1662_D));
  generic_pmos I_1631(.D(I_1695_D), .G(I_1631_G), .S(VDD));
  generic_nmos I_1632(.D(VSS), .G(I_1729_D), .S(I_1731_S));
  generic_pmos I_1633(.D(VDD), .G(I_1729_D), .S(I_1731_S));
  generic_nmos I_1634(.D(VSS), .G(I_1731_D), .S(I_1667_D));
  generic_pmos I_1635(.D(VDD), .G(I_1731_D), .S(I_1667_D));
  generic_nmos I_1636(.D(VSS), .G(I_1347_D), .S(I_1668_D));
  generic_pmos I_1637(.D(VDD), .G(I_1347_D), .S(I_1735_S));
  generic_nmos I_1638(.D(I_1638_D), .G(I_1347_D), .S(VSS));
  generic_pmos I_1639(.D(I_1733_S), .G(I_1347_D), .S(VDD));
  generic_nmos I_164(.D(I_261_D), .G(I_1187_S), .S(I_196_D));
  generic_nmos I_1640(.D(VSS), .G(I_1249_D), .S(I_1672_D));
  generic_pmos I_1641(.D(VDD), .G(I_1249_D), .S(I_1673_D));
  generic_nmos I_1642(.D(I_1642_D), .G(I_1643_G), .S(I_1674_D));
  generic_pmos I_1643(.D(I_1643_D), .G(I_1643_G), .S(I_1675_D));
  generic_nmos I_1644(.D(I_1644_D), .G(I_1645_G), .S(I_1676_D));
  generic_pmos I_1645(.D(I_1645_D), .G(I_1645_G), .S(I_1677_D));
  generic_nmos I_1646(.D(VSS), .G(I_1743_D), .S(I_1678_D));
  generic_pmos I_1647(.D(VDD), .G(I_1743_D), .S(I_1679_D));
  generic_nmos I_1648(.D(I_1648_D), .G(I_1679_D), .S(VSS));
  generic_pmos I_1649(.D(I_1649_D), .G(I_1679_D), .S(VDD));
  generic_pmos I_165(.D(VDD), .G(I_1187_S), .S(I_261_D));
  generic_nmos I_1650(.D(I_1650_D), .G(I_1651_G), .S(I_1682_D));
  generic_pmos I_1651(.D(I_1651_D), .G(I_1651_G), .S(I_1683_D));
  generic_nmos I_1652(.D(VSS), .G(I_151_D), .S(I_1685_D));
  generic_pmos I_1653(.D(VDD), .G(I_151_D), .S(I_1685_D));
  generic_nmos I_1654(.D(VSS), .G(I_151_D), .S(VSS));
  generic_pmos I_1655(.D(VDD), .G(I_151_D), .S(VDD));
  generic_nmos I_1656(.D(VSS), .G(I_1879_D), .S(I_1689_D));
  generic_pmos I_1657(.D(VDD), .G(I_1879_D), .S(I_1689_D));
  generic_nmos I_1658(.D(VSS), .G(I_1627_D), .S(I_1755_D));
  generic_pmos I_1659(.D(VDD), .G(I_1627_D), .S(I_1755_D));
  generic_nmos I_166(.D(I_263_D), .G(I_293_S), .S(VSS));
  generic_nmos I_1660(.D(I_1660_D), .G(I_1695_D), .S(I_1692_D));
  generic_pmos I_1661(.D(VDD), .G(I_1695_D), .S(I_1693_D));
  generic_nmos I_1662(.D(I_1662_D), .G(I_1598_S), .S(I_1694_D));
  generic_pmos I_1663(.D(VDD), .G(I_1598_S), .S(I_1695_D));
  generic_nmos I_1664(.D(I_1731_S), .G(I_1729_D), .S(VSS));
  generic_pmos I_1665(.D(I_1731_S), .G(I_1729_D), .S(VDD));
  generic_nmos I_1666(.D(I_1667_D), .G(I_1731_D), .S(VSS));
  generic_pmos I_1667(.D(I_1667_D), .G(I_1731_D), .S(VDD));
  generic_nmos I_1668(.D(I_1668_D), .G(I_1733_D), .S(I_1735_S));
  generic_pmos I_1669(.D(I_1735_S), .G(I_1733_D), .S(VDD));
  generic_pmos I_167(.D(I_263_D), .G(I_293_S), .S(VDD));
  generic_nmos I_1670(.D(VSS), .G(I_1735_D), .S(I_1671_S));
  generic_pmos I_1671(.D(VDD), .G(I_1735_D), .S(I_1671_S));
  generic_nmos I_1672(.D(I_1672_D), .G(I_1515_S), .S(I_1673_D));
  generic_pmos I_1673(.D(I_1673_D), .G(I_1515_S), .S(VDD));
  generic_nmos I_1674(.D(I_1674_D), .G(I_1675_G), .S(I_1674_S));
  generic_pmos I_1675(.D(I_1675_D), .G(I_1675_G), .S(I_1675_S));
  generic_nmos I_1676(.D(I_1676_D), .G(I_1677_G), .S(I_1676_S));
  generic_pmos I_1677(.D(I_1677_D), .G(I_1677_G), .S(I_1677_S));
  generic_nmos I_1678(.D(I_1678_D), .G(I_1807_D), .S(I_1679_D));
  generic_pmos I_1679(.D(I_1679_D), .G(I_1807_D), .S(VDD));
  generic_nmos I_168(.D(I_168_D), .G(I_169_G), .S(I_200_D));
  generic_nmos I_1680(.D(VSS), .G(I_1648_D), .S(I_1681_S));
  generic_pmos I_1681(.D(VDD), .G(I_1648_D), .S(I_1681_S));
  generic_nmos I_1682(.D(I_1682_D), .G(I_1683_G), .S(I_1682_S));
  generic_pmos I_1683(.D(I_1683_D), .G(I_1683_G), .S(I_1683_S));
  generic_nmos I_1684(.D(I_1685_D), .G(I_1685_G), .S(I_1684_S));
  generic_pmos I_1685(.D(I_1685_D), .G(I_1685_G), .S(I_1685_S));
  generic_nmos I_1686(.D(VSS), .G(I_1685_D), .S(I_1687_S));
  generic_pmos I_1687(.D(VDD), .G(I_1685_D), .S(I_1687_S));
  generic_nmos I_1688(.D(I_1689_D), .G(I_1879_D), .S(VSS));
  generic_pmos I_1689(.D(I_1689_D), .G(I_1879_D), .S(VDD));
  generic_pmos I_169(.D(I_169_D), .G(I_169_G), .S(I_201_D));
  generic_nmos I_1690(.D(I_1755_D), .G(I_1627_D), .S(VSS));
  generic_pmos I_1691(.D(I_1755_D), .G(I_1627_D), .S(VDD));
  generic_nmos I_1692(.D(I_1692_D), .G(I_1855_D), .S(VSS));
  generic_pmos I_1693(.D(I_1693_D), .G(I_1855_D), .S(VDD));
  generic_nmos I_1694(.D(I_1694_D), .G(I_1759_S), .S(VSS));
  generic_pmos I_1695(.D(I_1695_D), .G(I_1759_S), .S(VDD));
  generic_nmos I_1696(.D(I_1697_D), .G(I_1730_G), .S(I_1729_D));
  generic_pmos I_1697(.D(I_1697_D), .G(I_1761_D), .S(I_1729_D));
  generic_nmos I_1698(.D(I_1699_D), .G(I_1761_D), .S(I_1731_D));
  generic_pmos I_1699(.D(I_1699_D), .G(I_1730_G), .S(I_1731_D));
  generic_pmos I_17(.D(I_17_D), .G(I_17_G), .S(I_49_D));
  generic_nmos I_170(.D(I_235_D), .G(I_458_S), .S(I_202_D));
  generic_nmos I_1700(.D(I_1701_D), .G(I_1573_S), .S(I_1733_D));
  generic_pmos I_1701(.D(I_1701_D), .G(I_1511_S), .S(I_1733_D));
  generic_nmos I_1702(.D(I_1733_S), .G(I_1511_S), .S(I_1735_D));
  generic_pmos I_1703(.D(I_1733_S), .G(I_1573_S), .S(I_1735_D));
  generic_nmos I_1704(.D(VSS), .G(I_1609_D), .S(I_1736_D));
  generic_pmos I_1705(.D(VDD), .G(I_1515_S), .S(I_1737_D));
  generic_nmos I_1706(.D(I_1706_D), .G(I_1706_G), .S(I_1738_D));
  generic_pmos I_1707(.D(I_1707_D), .G(I_1738_G), .S(I_1739_D));
  generic_nmos I_1708(.D(I_1741_S), .G(I_3013_S), .S(VSS));
  generic_pmos I_1709(.D(I_1709_D), .G(I_1740_G), .S(VDD));
  generic_pmos I_171(.D(I_235_D), .G(I_458_S), .S(VDD));
  generic_nmos I_1710(.D(I_1743_D), .G(I_1839_S), .S(I_1742_D));
  generic_pmos I_1711(.D(VDD), .G(I_1741_S), .S(I_1743_D));
  generic_nmos I_1712(.D(VSS), .G(I_1648_D), .S(I_2545_S));
  generic_pmos I_1713(.D(I_1713_D), .G(I_1744_G), .S(I_2545_S));
  generic_nmos I_1714(.D(VSS), .G(I_2133_G), .S(VSS));
  generic_pmos I_1715(.D(I_1715_D), .G(I_1746_G), .S(VDD));
  generic_nmos I_1716(.D(I_1749_S), .G(I_1748_S), .S(VSS));
  generic_pmos I_1717(.D(I_1748_S), .G(I_1751_S), .S(VDD));
  generic_nmos I_1718(.D(I_1751_S), .G(I_1750_S), .S(VSS));
  generic_pmos I_1719(.D(I_1750_S), .G(I_151_D), .S(VDD));
  generic_nmos I_172(.D(I_172_D), .G(I_173_G), .S(I_204_D));
  generic_nmos I_1720(.D(I_1753_S), .G(I_1752_S), .S(VSS));
  generic_pmos I_1721(.D(I_1752_S), .G(I_1751_S), .S(VDD));
  generic_nmos I_1722(.D(VSS), .G(I_1627_D), .S(I_1755_D));
  generic_pmos I_1723(.D(VDD), .G(I_1627_D), .S(I_1755_D));
  generic_nmos I_1724(.D(VSS), .G(I_1915_S), .S(I_1757_D));
  generic_pmos I_1725(.D(VDD), .G(I_1915_S), .S(I_1757_D));
  generic_nmos I_1726(.D(I_1759_S), .G(I_1758_S), .S(VSS));
  generic_pmos I_1727(.D(I_1758_S), .G(I_1821_D), .S(VDD));
  generic_nmos I_1728(.D(I_1729_D), .G(I_1761_D), .S(I_1729_S));
  generic_pmos I_1729(.D(I_1729_D), .G(I_1730_G), .S(I_1729_S));
  generic_pmos I_173(.D(I_173_D), .G(I_173_G), .S(I_205_D));
  generic_nmos I_1730(.D(I_1731_D), .G(I_1730_G), .S(I_1731_S));
  generic_pmos I_1731(.D(I_1731_D), .G(I_1761_D), .S(I_1731_S));
  generic_nmos I_1732(.D(I_1733_D), .G(I_1511_S), .S(I_1733_S));
  generic_pmos I_1733(.D(I_1733_D), .G(I_1573_S), .S(I_1733_S));
  generic_nmos I_1734(.D(I_1735_D), .G(I_1573_S), .S(I_1735_S));
  generic_pmos I_1735(.D(I_1735_D), .G(I_1511_S), .S(I_1735_S));
  generic_nmos I_1736(.D(I_1736_D), .G(I_1515_S), .S(I_1737_D));
  generic_pmos I_1737(.D(I_1737_D), .G(I_1609_D), .S(VDD));
  generic_nmos I_1738(.D(I_1738_D), .G(I_1738_G), .S(I_1738_S));
  generic_pmos I_1739(.D(I_1739_D), .G(I_1739_G), .S(I_1739_S));
  generic_nmos I_174(.D(I_174_D), .G(I_175_G), .S(I_206_D));
  generic_nmos I_1740(.D(VSS), .G(I_1740_G), .S(I_1740_S));
  generic_pmos I_1741(.D(VDD), .G(I_3013_S), .S(I_1741_S));
  generic_nmos I_1742(.D(I_1742_D), .G(I_1741_S), .S(VSS));
  generic_pmos I_1743(.D(I_1743_D), .G(I_1839_S), .S(VDD));
  generic_nmos I_1744(.D(I_2545_S), .G(I_1744_G), .S(I_1744_S));
  generic_pmos I_1745(.D(I_2545_S), .G(I_1585_D), .S(VDD));
  generic_nmos I_1746(.D(VSS), .G(I_1746_G), .S(I_1746_S));
  generic_pmos I_1747(.D(VDD), .G(I_2133_G), .S(VDD));
  generic_nmos I_1748(.D(VSS), .G(I_1751_S), .S(I_1748_S));
  generic_pmos I_1749(.D(VDD), .G(I_1748_S), .S(I_1749_S));
  generic_pmos I_175(.D(I_175_D), .G(I_175_G), .S(I_207_D));
  generic_nmos I_1750(.D(VSS), .G(I_151_D), .S(I_1750_S));
  generic_pmos I_1751(.D(VDD), .G(I_1750_S), .S(I_1751_S));
  generic_nmos I_1752(.D(VSS), .G(I_1751_S), .S(I_1752_S));
  generic_pmos I_1753(.D(VDD), .G(I_1752_S), .S(I_1753_S));
  generic_nmos I_1754(.D(I_1755_D), .G(I_1627_D), .S(VSS));
  generic_pmos I_1755(.D(I_1755_D), .G(I_1627_D), .S(VDD));
  generic_nmos I_1756(.D(I_1757_D), .G(I_1915_S), .S(VSS));
  generic_pmos I_1757(.D(I_1757_D), .G(I_1915_S), .S(VDD));
  generic_nmos I_1758(.D(VSS), .G(I_1821_D), .S(I_1758_S));
  generic_pmos I_1759(.D(VDD), .G(I_1758_S), .S(I_1759_S));
  generic_nmos I_176(.D(I_176_D), .G(I_177_G), .S(I_208_D));
  generic_nmos I_1760(.D(I_1761_D), .G(I_1761_G), .S(VSS));
  generic_pmos I_1761(.D(I_1761_D), .G(I_1761_G), .S(VDD));
  generic_nmos I_1762(.D(I_1763_D), .G(I_1831_S), .S(VSS));
  generic_pmos I_1763(.D(I_1763_D), .G(I_1831_S), .S(VDD));
  generic_nmos I_1764(.D(I_1861_D), .G(I_1895_S), .S(VSS));
  generic_pmos I_1765(.D(I_1861_D), .G(I_1895_S), .S(VDD));
  generic_nmos I_1766(.D(I_1893_S), .G(I_1831_S), .S(I_1798_D));
  generic_pmos I_1767(.D(VDD), .G(I_1831_S), .S(I_1893_S));
  generic_nmos I_1768(.D(VSS), .G(I_1673_D), .S(I_1800_D));
  generic_pmos I_1769(.D(VDD), .G(I_1673_D), .S(I_1832_D));
  generic_pmos I_177(.D(I_177_D), .G(I_177_G), .S(I_209_D));
  generic_nmos I_1770(.D(I_1770_D), .G(I_1771_G), .S(I_1802_D));
  generic_pmos I_1771(.D(I_1771_D), .G(I_1771_G), .S(I_1803_D));
  generic_nmos I_1772(.D(I_1772_D), .G(I_1773_G), .S(I_1804_D));
  generic_pmos I_1773(.D(I_1773_D), .G(I_1773_G), .S(I_1805_D));
  generic_nmos I_1774(.D(I_1807_D), .G(I_3431_S), .S(I_1806_D));
  generic_pmos I_1775(.D(VDD), .G(I_3431_S), .S(I_1807_D));
  generic_nmos I_1776(.D(I_2065_S), .G(I_1681_S), .S(I_1808_D));
  generic_pmos I_1777(.D(VDD), .G(I_1681_S), .S(I_2065_S));
  generic_nmos I_1778(.D(I_1778_D), .G(I_1779_G), .S(I_1810_D));
  generic_pmos I_1779(.D(I_1779_D), .G(I_1779_G), .S(I_1811_D));
  generic_nmos I_178(.D(I_178_D), .G(I_179_G), .S(I_210_D));
  generic_nmos I_1780(.D(I_1845_D), .G(I_1051_S), .S(I_1812_D));
  generic_pmos I_1781(.D(I_1845_D), .G(I_1051_S), .S(VDD));
  generic_nmos I_1782(.D(I_1879_D), .G(I_1847_D), .S(VSS));
  generic_pmos I_1783(.D(I_1879_D), .G(I_1847_D), .S(VDD));
  generic_nmos I_1784(.D(I_1881_D), .G(I_1911_S), .S(VSS));
  generic_pmos I_1785(.D(I_1881_D), .G(I_1911_S), .S(VDD));
  generic_nmos I_1786(.D(VSS), .G(I_1853_S), .S(I_1821_D));
  generic_pmos I_1787(.D(VDD), .G(I_1853_S), .S(I_1821_D));
  generic_nmos I_1788(.D(VSS), .G(I_1853_S), .S(I_1821_D));
  generic_pmos I_1789(.D(VDD), .G(I_1853_S), .S(I_1821_D));
  generic_pmos I_179(.D(I_179_D), .G(I_179_G), .S(I_211_D));
  generic_nmos I_1790(.D(I_1855_D), .G(I_1599_S), .S(I_1822_D));
  generic_pmos I_1791(.D(I_1855_D), .G(I_1599_S), .S(VDD));
  generic_nmos I_1792(.D(VSS), .G(I_1345_D), .S(I_1825_D));
  generic_pmos I_1793(.D(VDD), .G(I_1345_D), .S(I_1825_D));
  generic_nmos I_1794(.D(VSS), .G(I_1763_D), .S(I_1826_D));
  generic_pmos I_1795(.D(VDD), .G(I_1763_D), .S(I_1891_S));
  generic_nmos I_1796(.D(VSS), .G(I_1347_D), .S(I_1828_D));
  generic_pmos I_1797(.D(VDD), .G(I_1347_D), .S(I_1895_S));
  generic_nmos I_1798(.D(I_1798_D), .G(I_1347_D), .S(VSS));
  generic_pmos I_1799(.D(I_1893_S), .G(I_1347_D), .S(VDD));
  generic_nmos I_18(.D(I_18_D), .G(I_19_G), .S(I_50_D));
  generic_nmos I_180(.D(I_245_D), .G(I_277_D), .S(VSS));
  generic_nmos I_1800(.D(I_1800_D), .G(I_1737_D), .S(I_1832_D));
  generic_pmos I_1801(.D(I_1832_D), .G(I_1737_D), .S(VDD));
  generic_nmos I_1802(.D(I_1802_D), .G(I_1803_G), .S(I_1834_D));
  generic_pmos I_1803(.D(I_1803_D), .G(I_1803_G), .S(I_1835_D));
  generic_nmos I_1804(.D(I_1804_D), .G(I_1805_G), .S(I_1836_D));
  generic_pmos I_1805(.D(I_1805_D), .G(I_1805_G), .S(I_1837_D));
  generic_nmos I_1806(.D(I_1806_D), .G(I_2253_D), .S(VSS));
  generic_pmos I_1807(.D(I_1807_D), .G(I_2253_D), .S(VDD));
  generic_nmos I_1808(.D(I_1808_D), .G(I_1585_D), .S(VSS));
  generic_pmos I_1809(.D(I_2065_S), .G(I_1585_D), .S(VDD));
  generic_pmos I_181(.D(I_245_D), .G(I_277_D), .S(VDD));
  generic_nmos I_1810(.D(I_1810_D), .G(I_1811_G), .S(VSS));
  generic_pmos I_1811(.D(I_1811_D), .G(I_1811_G), .S(VDD));
  generic_nmos I_1812(.D(I_1812_D), .G(I_1397_D), .S(I_1844_D));
  generic_pmos I_1813(.D(VDD), .G(I_1397_D), .S(I_1845_D));
  generic_nmos I_1814(.D(VSS), .G(I_1911_D), .S(I_1847_D));
  generic_pmos I_1815(.D(VDD), .G(I_1911_D), .S(I_1847_D));
  generic_nmos I_1816(.D(VSS), .G(I_1913_D), .S(I_1911_S));
  generic_pmos I_1817(.D(VDD), .G(I_1913_D), .S(I_1911_S));
  generic_nmos I_1818(.D(I_1821_D), .G(I_1853_S), .S(VSS));
  generic_pmos I_1819(.D(I_1821_D), .G(I_1853_S), .S(VDD));
  generic_nmos I_182(.D(I_279_D), .G(I_247_D), .S(VSS));
  generic_nmos I_1820(.D(I_1821_D), .G(I_1853_S), .S(VSS));
  generic_pmos I_1821(.D(I_1821_D), .G(I_1853_S), .S(VDD));
  generic_nmos I_1822(.D(I_1822_D), .G(I_1758_S), .S(I_1854_D));
  generic_pmos I_1823(.D(VDD), .G(I_1758_S), .S(I_1855_D));
  generic_nmos I_1824(.D(I_1825_D), .G(I_1345_D), .S(VSS));
  generic_pmos I_1825(.D(I_1825_D), .G(I_1345_D), .S(VDD));
  generic_nmos I_1826(.D(I_1826_D), .G(I_2311_S), .S(I_1858_D));
  generic_pmos I_1827(.D(I_1891_S), .G(I_2311_S), .S(VDD));
  generic_nmos I_1828(.D(I_1828_D), .G(I_1893_D), .S(I_1895_S));
  generic_pmos I_1829(.D(I_1895_S), .G(I_1893_D), .S(VDD));
  generic_pmos I_183(.D(I_279_D), .G(I_247_D), .S(VDD));
  generic_nmos I_1830(.D(VSS), .G(I_1895_D), .S(I_1831_S));
  generic_pmos I_1831(.D(VDD), .G(I_1895_D), .S(I_1831_S));
  generic_nmos I_1832(.D(I_1832_D), .G(I_1833_G), .S(I_1832_S));
  generic_pmos I_1833(.D(VDD), .G(I_1833_G), .S(I_1833_S));
  generic_nmos I_1834(.D(I_1834_D), .G(I_1835_G), .S(I_1834_S));
  generic_pmos I_1835(.D(I_1835_D), .G(I_1835_G), .S(I_1835_S));
  generic_nmos I_1836(.D(I_1836_D), .G(I_1837_G), .S(I_1836_S));
  generic_pmos I_1837(.D(I_1837_D), .G(I_1837_G), .S(I_1837_S));
  generic_nmos I_1838(.D(VSS), .G(I_2253_D), .S(I_1839_S));
  generic_pmos I_1839(.D(VDD), .G(I_2253_D), .S(I_1839_S));
  generic_nmos I_184(.D(I_185_D), .G(I_281_D), .S(VSS));
  generic_nmos I_1840(.D(VSS), .G(I_2065_S), .S(I_2033_D));
  generic_pmos I_1841(.D(VDD), .G(I_2065_S), .S(I_2033_D));
  generic_nmos I_1842(.D(VSS), .G(I_1425_S), .S(I_1843_S));
  generic_pmos I_1843(.D(VDD), .G(I_1425_S), .S(I_1843_S));
  generic_nmos I_1844(.D(I_1844_D), .G(I_457_D), .S(VSS));
  generic_pmos I_1845(.D(I_1845_D), .G(I_457_D), .S(VDD));
  generic_nmos I_1846(.D(I_1847_D), .G(I_1911_D), .S(VSS));
  generic_pmos I_1847(.D(I_1847_D), .G(I_1911_D), .S(VDD));
  generic_nmos I_1848(.D(I_1911_S), .G(I_1913_D), .S(VSS));
  generic_pmos I_1849(.D(I_1911_S), .G(I_1913_D), .S(VDD));
  generic_pmos I_185(.D(I_185_D), .G(I_281_D), .S(VDD));
  generic_nmos I_1850(.D(VSS), .G(I_1279_S), .S(I_1853_S));
  generic_pmos I_1851(.D(VDD), .G(I_1279_S), .S(I_1853_S));
  generic_nmos I_1852(.D(VSS), .G(I_1279_S), .S(I_1853_S));
  generic_pmos I_1853(.D(VDD), .G(I_1279_S), .S(I_1853_S));
  generic_nmos I_1854(.D(I_1854_D), .G(I_1901_D), .S(VSS));
  generic_pmos I_1855(.D(I_1855_D), .G(I_1901_D), .S(VDD));
  generic_nmos I_1856(.D(I_1889_D), .G(I_1987_D), .S(I_1888_D));
  generic_pmos I_1857(.D(VDD), .G(I_1888_G), .S(I_1889_D));
  generic_nmos I_1858(.D(I_1858_D), .G(I_1923_D), .S(I_1890_D));
  generic_pmos I_1859(.D(I_1891_S), .G(I_2151_S), .S(VDD));
  generic_nmos I_186(.D(VSS), .G(I_347_D), .S(I_251_S));
  generic_nmos I_1860(.D(I_1861_D), .G(I_1733_S), .S(I_1893_D));
  generic_pmos I_1861(.D(I_1861_D), .G(I_1671_S), .S(I_1893_D));
  generic_nmos I_1862(.D(I_1893_S), .G(I_1671_S), .S(I_1895_D));
  generic_pmos I_1863(.D(I_1893_S), .G(I_1733_S), .S(I_1895_D));
  generic_nmos I_1864(.D(I_1864_D), .G(I_1864_G), .S(I_1896_D));
  generic_pmos I_1865(.D(I_1865_D), .G(I_1896_G), .S(I_1897_D));
  generic_nmos I_1866(.D(VSS), .G(I_873_D), .S(I_1899_S));
  generic_pmos I_1867(.D(VDD), .G(I_101_D), .S(I_1899_D));
  generic_nmos I_1868(.D(I_1901_D), .G(I_2157_S), .S(I_1900_D));
  generic_pmos I_1869(.D(VDD), .G(I_101_D), .S(I_1901_D));
  generic_pmos I_187(.D(VDD), .G(I_347_D), .S(I_251_S));
  generic_nmos I_1870(.D(I_1870_D), .G(I_1870_G), .S(I_1902_D));
  generic_pmos I_1871(.D(I_1871_D), .G(I_1902_G), .S(I_1903_D));
  generic_nmos I_1872(.D(I_2545_S), .G(I_2033_D), .S(I_1906_S));
  generic_pmos I_1873(.D(I_1873_D), .G(I_1904_G), .S(I_2545_S));
  generic_nmos I_1874(.D(I_1874_D), .G(I_1874_G), .S(VSS));
  generic_pmos I_1875(.D(I_1906_S), .G(I_1843_S), .S(VDD));
  generic_nmos I_1876(.D(I_1876_D), .G(I_1876_G), .S(VSS));
  generic_pmos I_1877(.D(I_1908_S), .G(I_503_D), .S(VDD));
  generic_nmos I_1878(.D(I_1879_D), .G(I_1908_S), .S(I_1911_D));
  generic_pmos I_1879(.D(I_1879_D), .G(I_503_D), .S(I_1911_D));
  generic_nmos I_188(.D(I_285_D), .G(I_157_D), .S(I_220_D));
  generic_nmos I_1880(.D(I_1881_D), .G(I_503_D), .S(I_1913_D));
  generic_pmos I_1881(.D(I_1881_D), .G(I_1908_S), .S(I_1913_D));
  generic_nmos I_1882(.D(VSS), .G(I_1853_S), .S(I_1915_S));
  generic_pmos I_1883(.D(VDD), .G(I_1879_D), .S(I_1915_D));
  generic_nmos I_1884(.D(VSS), .G(I_1949_D), .S(I_1916_D));
  generic_pmos I_1885(.D(VDD), .G(I_1693_D), .S(I_1917_D));
  generic_nmos I_1886(.D(VSS), .G(I_2077_D), .S(I_1919_D));
  generic_pmos I_1887(.D(VDD), .G(I_2077_D), .S(I_1919_D));
  generic_nmos I_1888(.D(I_1888_D), .G(I_1888_G), .S(VSS));
  generic_pmos I_1889(.D(I_1889_D), .G(I_1987_D), .S(VDD));
  generic_pmos I_189(.D(VDD), .G(I_157_D), .S(I_285_D));
  generic_nmos I_1890(.D(I_1890_D), .G(I_2151_S), .S(I_1891_S));
  generic_pmos I_1891(.D(VDD), .G(I_1923_D), .S(I_1891_S));
  generic_nmos I_1892(.D(I_1893_D), .G(I_1671_S), .S(I_1893_S));
  generic_pmos I_1893(.D(I_1893_D), .G(I_1733_S), .S(I_1893_S));
  generic_nmos I_1894(.D(I_1895_D), .G(I_1733_S), .S(I_1895_S));
  generic_pmos I_1895(.D(I_1895_D), .G(I_1671_S), .S(I_1895_S));
  generic_nmos I_1896(.D(I_1896_D), .G(I_1896_G), .S(I_1896_S));
  generic_pmos I_1897(.D(I_1897_D), .G(I_1897_G), .S(I_1897_S));
  generic_nmos I_1898(.D(I_1899_S), .G(I_101_D), .S(VSS));
  generic_pmos I_1899(.D(I_1899_D), .G(I_873_D), .S(I_1899_S));
  generic_pmos I_19(.D(I_19_D), .G(I_19_G), .S(I_51_D));
  generic_nmos I_190(.D(I_190_D), .G(I_191_G), .S(I_222_D));
  generic_nmos I_1900(.D(I_1900_D), .G(I_101_D), .S(VSS));
  generic_pmos I_1901(.D(I_1901_D), .G(I_2157_S), .S(VDD));
  generic_nmos I_1902(.D(I_1902_D), .G(I_1902_G), .S(I_1902_S));
  generic_pmos I_1903(.D(I_1903_D), .G(I_1903_G), .S(I_1903_S));
  generic_nmos I_1904(.D(I_1906_S), .G(I_1904_G), .S(I_1904_S));
  generic_pmos I_1905(.D(I_2545_S), .G(I_2065_S), .S(I_1906_S));
  generic_nmos I_1906(.D(VSS), .G(I_1843_S), .S(I_1906_S));
  generic_pmos I_1907(.D(VDD), .G(I_1907_G), .S(I_1907_S));
  generic_nmos I_1908(.D(VSS), .G(I_503_D), .S(I_1908_S));
  generic_pmos I_1909(.D(VDD), .G(I_1909_G), .S(I_1909_S));
  generic_pmos I_191(.D(I_191_D), .G(I_191_G), .S(I_223_D));
  generic_nmos I_1910(.D(I_1911_D), .G(I_503_D), .S(I_1911_S));
  generic_pmos I_1911(.D(I_1911_D), .G(I_1908_S), .S(I_1911_S));
  generic_nmos I_1912(.D(I_1913_D), .G(I_1908_S), .S(I_1913_S));
  generic_pmos I_1913(.D(I_1913_D), .G(I_503_D), .S(I_1913_S));
  generic_nmos I_1914(.D(I_1915_S), .G(I_1879_D), .S(VSS));
  generic_pmos I_1915(.D(I_1915_D), .G(I_1853_S), .S(I_1915_S));
  generic_nmos I_1916(.D(I_1916_D), .G(I_1693_D), .S(I_1917_D));
  generic_pmos I_1917(.D(I_1917_D), .G(I_1949_D), .S(VDD));
  generic_nmos I_1918(.D(I_1919_D), .G(I_2077_D), .S(VSS));
  generic_pmos I_1919(.D(I_1919_D), .G(I_2077_D), .S(VDD));
  generic_nmos I_192(.D(I_225_D), .G(I_227_D), .S(I_224_D));
  generic_nmos I_1920(.D(I_2209_S), .G(I_1921_G), .S(I_1952_D));
  generic_pmos I_1921(.D(VDD), .G(I_1921_G), .S(I_2209_S));
  generic_nmos I_1922(.D(I_1923_D), .G(I_1991_S), .S(VSS));
  generic_pmos I_1923(.D(I_1923_D), .G(I_1991_S), .S(VDD));
  generic_nmos I_1924(.D(I_2021_D), .G(I_2055_S), .S(VSS));
  generic_pmos I_1925(.D(I_2021_D), .G(I_2055_S), .S(VDD));
  generic_nmos I_1926(.D(I_2053_S), .G(I_1991_S), .S(I_1958_D));
  generic_pmos I_1927(.D(VDD), .G(I_1991_S), .S(I_2053_S));
  generic_nmos I_1928(.D(I_1928_D), .G(I_1929_G), .S(I_1960_D));
  generic_pmos I_1929(.D(I_1929_D), .G(I_1929_G), .S(I_1961_D));
  generic_pmos I_193(.D(I_193_D), .G(I_227_D), .S(I_225_D));
  generic_nmos I_1930(.D(VSS), .G(I_1899_S), .S(I_1962_D));
  generic_pmos I_1931(.D(I_1962_D), .G(I_1899_S), .S(I_1995_S));
  generic_nmos I_1932(.D(I_1997_D), .G(I_2317_S), .S(VSS));
  generic_pmos I_1933(.D(I_1997_D), .G(I_2317_S), .S(VDD));
  generic_nmos I_1934(.D(I_1934_D), .G(I_1935_G), .S(VSS));
  generic_pmos I_1935(.D(I_1935_D), .G(I_1935_G), .S(VDD));
  generic_nmos I_1936(.D(I_1936_D), .G(I_1937_G), .S(I_1969_D));
  generic_pmos I_1937(.D(I_1937_D), .G(I_1937_G), .S(I_1969_D));
  generic_nmos I_1938(.D(I_1938_D), .G(I_1939_G), .S(I_1970_D));
  generic_pmos I_1939(.D(I_1939_D), .G(I_1939_G), .S(I_1971_D));
  generic_nmos I_194(.D(VSS), .G(I_291_D), .S(I_226_D));
  generic_nmos I_1940(.D(VSS), .G(I_1943_D), .S(I_1973_D));
  generic_pmos I_1941(.D(VDD), .G(I_1943_D), .S(I_1973_D));
  generic_nmos I_1942(.D(I_1943_D), .G(I_1309_D), .S(VSS));
  generic_pmos I_1943(.D(I_1943_D), .G(I_1309_D), .S(VDD));
  generic_nmos I_1944(.D(I_2009_D), .G(I_1879_D), .S(VSS));
  generic_pmos I_1945(.D(I_2009_D), .G(I_1879_D), .S(VDD));
  generic_nmos I_1946(.D(I_1946_D), .G(I_1947_G), .S(VSS));
  generic_pmos I_1947(.D(I_1947_D), .G(I_1947_G), .S(VDD));
  generic_nmos I_1948(.D(I_1949_D), .G(I_1689_D), .S(VSS));
  generic_pmos I_1949(.D(I_1949_D), .G(I_1689_D), .S(VDD));
  generic_pmos I_195(.D(VDD), .G(I_291_D), .S(I_227_D));
  generic_nmos I_1950(.D(I_2015_D), .G(I_3669_D), .S(I_1982_D));
  generic_pmos I_1951(.D(I_2015_D), .G(I_3669_D), .S(VDD));
  generic_nmos I_1952(.D(I_1952_D), .G(I_1985_S), .S(VSS));
  generic_pmos I_1953(.D(I_2209_S), .G(I_1985_S), .S(VDD));
  generic_nmos I_1954(.D(VSS), .G(I_2051_D), .S(I_1986_D));
  generic_pmos I_1955(.D(VDD), .G(I_2051_D), .S(I_1987_D));
  generic_nmos I_1956(.D(VSS), .G(I_1347_D), .S(I_1988_D));
  generic_pmos I_1957(.D(VDD), .G(I_1347_D), .S(I_2055_S));
  generic_nmos I_1958(.D(I_1958_D), .G(I_1347_D), .S(VSS));
  generic_pmos I_1959(.D(I_2053_S), .G(I_1347_D), .S(VDD));
  generic_nmos I_196(.D(I_196_D), .G(I_229_S), .S(VSS));
  generic_nmos I_1960(.D(I_1960_D), .G(I_1961_G), .S(I_1992_D));
  generic_pmos I_1961(.D(I_1961_D), .G(I_1961_G), .S(I_1993_D));
  generic_nmos I_1962(.D(I_1962_D), .G(I_101_D), .S(I_1994_D));
  generic_pmos I_1963(.D(I_1995_S), .G(I_101_D), .S(VDD));
  generic_nmos I_1964(.D(VSS), .G(I_2317_S), .S(I_1997_D));
  generic_pmos I_1965(.D(VDD), .G(I_2317_S), .S(I_1997_D));
  generic_nmos I_1966(.D(VSS), .G(I_2063_D), .S(I_1998_D));
  generic_pmos I_1967(.D(VDD), .G(I_2063_D), .S(I_1999_D));
  generic_nmos I_1968(.D(I_1969_D), .G(I_1906_S), .S(VSS));
  generic_pmos I_1969(.D(I_1969_D), .G(I_1906_S), .S(VDD));
  generic_pmos I_197(.D(I_261_D), .G(I_229_S), .S(VDD));
  generic_nmos I_1970(.D(I_1970_D), .G(I_1971_G), .S(I_2002_D));
  generic_pmos I_1971(.D(I_1971_D), .G(I_1971_G), .S(I_2003_D));
  generic_nmos I_1972(.D(I_1973_D), .G(I_1943_D), .S(VSS));
  generic_pmos I_1973(.D(I_1973_D), .G(I_1943_D), .S(VDD));
  generic_nmos I_1974(.D(VSS), .G(I_1973_D), .S(I_2007_D));
  generic_pmos I_1975(.D(VDD), .G(I_1973_D), .S(I_2007_D));
  generic_nmos I_1976(.D(VSS), .G(I_1879_D), .S(I_2009_D));
  generic_pmos I_1977(.D(VDD), .G(I_1879_D), .S(I_2009_D));
  generic_nmos I_1978(.D(VSS), .G(I_2075_D), .S(I_2010_D));
  generic_pmos I_1979(.D(VDD), .G(I_2075_D), .S(I_2011_D));
  generic_nmos I_198(.D(VSS), .G(I_1187_S), .S(I_230_D));
  generic_nmos I_1980(.D(VSS), .G(I_1689_D), .S(I_2012_D));
  generic_pmos I_1981(.D(VDD), .G(I_1689_D), .S(I_2013_D));
  generic_nmos I_1982(.D(I_1982_D), .G(I_2238_S), .S(I_2014_D));
  generic_pmos I_1983(.D(VDD), .G(I_2238_S), .S(I_2015_D));
  generic_nmos I_1984(.D(VSS), .G(I_2049_D), .S(I_1985_S));
  generic_pmos I_1985(.D(VDD), .G(I_2049_D), .S(I_1985_S));
  generic_nmos I_1986(.D(I_1986_D), .G(I_2115_D), .S(I_1987_D));
  generic_pmos I_1987(.D(I_1987_D), .G(I_2115_D), .S(VDD));
  generic_nmos I_1988(.D(I_1988_D), .G(I_2053_D), .S(I_2055_S));
  generic_pmos I_1989(.D(I_2055_S), .G(I_2053_D), .S(VDD));
  generic_pmos I_199(.D(VDD), .G(I_1187_S), .S(I_293_S));
  generic_nmos I_1990(.D(VSS), .G(I_2055_D), .S(I_1991_S));
  generic_pmos I_1991(.D(VDD), .G(I_2055_D), .S(I_1991_S));
  generic_nmos I_1992(.D(I_1992_D), .G(I_1993_G), .S(I_1992_S));
  generic_pmos I_1993(.D(I_1993_D), .G(I_1993_G), .S(I_1993_S));
  generic_nmos I_1994(.D(I_1994_D), .G(I_873_D), .S(VSS));
  generic_pmos I_1995(.D(VDD), .G(I_873_D), .S(I_1995_S));
  generic_nmos I_1996(.D(I_1997_D), .G(I_2317_S), .S(VSS));
  generic_pmos I_1997(.D(I_1997_D), .G(I_2317_S), .S(VDD));
  generic_nmos I_1998(.D(I_1998_D), .G(I_2127_D), .S(I_1999_D));
  generic_pmos I_1999(.D(I_1999_D), .G(I_2127_D), .S(VDD));
  generic_nmos I_2(.D(I_3_D), .G(I_3_G), .S(VSS));
  generic_nmos I_20(.D(I_20_D), .G(I_21_G), .S(I_52_D));
  generic_nmos I_200(.D(I_200_D), .G(I_201_G), .S(I_232_D));
  generic_nmos I_2000(.D(VSS), .G(I_1969_D), .S(I_2001_S));
  generic_pmos I_2001(.D(VDD), .G(I_1969_D), .S(I_2001_S));
  generic_nmos I_2002(.D(I_2002_D), .G(I_2003_G), .S(I_2002_S));
  generic_pmos I_2003(.D(I_2003_D), .G(I_2003_G), .S(I_2003_S));
  generic_nmos I_2004(.D(VSS), .G(I_2005_G), .S(I_2004_S));
  generic_pmos I_2005(.D(VDD), .G(I_2005_G), .S(I_2005_S));
  generic_nmos I_2006(.D(I_2007_D), .G(I_1973_D), .S(VSS));
  generic_pmos I_2007(.D(I_2007_D), .G(I_1973_D), .S(VDD));
  generic_nmos I_2008(.D(I_2009_D), .G(I_1879_D), .S(VSS));
  generic_pmos I_2009(.D(I_2009_D), .G(I_1879_D), .S(VDD));
  generic_pmos I_201(.D(I_201_D), .G(I_201_G), .S(I_233_D));
  generic_nmos I_2010(.D(I_2010_D), .G(I_2139_D), .S(I_2011_D));
  generic_pmos I_2011(.D(I_2011_D), .G(I_2139_D), .S(VDD));
  generic_nmos I_2012(.D(I_2012_D), .G(I_2011_D), .S(I_2013_D));
  generic_pmos I_2013(.D(I_2013_D), .G(I_2011_D), .S(VDD));
  generic_nmos I_2014(.D(I_2014_D), .G(I_2078_S), .S(VSS));
  generic_pmos I_2015(.D(I_2015_D), .G(I_2078_S), .S(VDD));
  generic_nmos I_2016(.D(I_2209_S), .G(I_2305_S), .S(I_2049_D));
  generic_pmos I_2017(.D(I_2209_S), .G(I_2529_S), .S(I_2049_D));
  generic_nmos I_2018(.D(I_2051_D), .G(I_2147_S), .S(I_2050_D));
  generic_pmos I_2019(.D(VDD), .G(I_2050_G), .S(I_2051_D));
  generic_nmos I_202(.D(I_202_D), .G(I_297_S), .S(I_234_D));
  generic_nmos I_2020(.D(I_2021_D), .G(I_1893_S), .S(I_2053_D));
  generic_pmos I_2021(.D(I_2021_D), .G(I_1831_S), .S(I_2053_D));
  generic_nmos I_2022(.D(I_2053_S), .G(I_1831_S), .S(I_2055_D));
  generic_pmos I_2023(.D(I_2053_S), .G(I_1893_S), .S(I_2055_D));
  generic_nmos I_2024(.D(I_2024_D), .G(I_2024_G), .S(I_2056_D));
  generic_pmos I_2025(.D(I_2025_D), .G(I_2056_G), .S(I_2057_D));
  generic_nmos I_2026(.D(I_2026_D), .G(I_2026_G), .S(VSS));
  generic_pmos I_2027(.D(I_2058_S), .G(I_2699_D), .S(VDD));
  generic_nmos I_2028(.D(I_2028_D), .G(I_2028_G), .S(I_2060_D));
  generic_pmos I_2029(.D(I_2029_D), .G(I_2060_G), .S(I_2061_D));
  generic_pmos I_203(.D(VDD), .G(I_297_S), .S(I_235_D));
  generic_nmos I_2030(.D(I_2063_D), .G(I_2159_S), .S(I_2062_D));
  generic_pmos I_2031(.D(VDD), .G(I_2062_G), .S(I_2063_D));
  generic_nmos I_2032(.D(I_2033_D), .G(I_1969_D), .S(I_2709_S));
  generic_pmos I_2033(.D(I_2033_D), .G(I_2001_S), .S(I_2709_S));
  generic_nmos I_2034(.D(I_2034_D), .G(I_2034_G), .S(I_2066_D));
  generic_pmos I_2035(.D(I_2035_D), .G(I_2066_G), .S(I_2067_D));
  generic_nmos I_2036(.D(I_2069_D), .G(I_1518_D), .S(I_2068_D));
  generic_pmos I_2037(.D(VDD), .G(I_2133_G), .S(I_2069_D));
  generic_nmos I_2038(.D(I_2167_S), .G(I_2231_D), .S(I_2071_D));
  generic_pmos I_2039(.D(I_2167_S), .G(I_2103_D), .S(I_2071_D));
  generic_nmos I_204(.D(I_204_D), .G(I_205_G), .S(I_236_D));
  generic_nmos I_2040(.D(I_2041_D), .G(I_1973_D), .S(I_2073_D));
  generic_pmos I_2041(.D(I_2041_D), .G(I_2007_D), .S(I_2073_D));
  generic_nmos I_2042(.D(I_2075_D), .G(I_2171_S), .S(I_2074_D));
  generic_pmos I_2043(.D(VDD), .G(I_2071_D), .S(I_2075_D));
  generic_nmos I_2044(.D(I_2077_D), .G(I_2013_D), .S(I_2076_D));
  generic_pmos I_2045(.D(VDD), .G(I_1917_D), .S(I_2077_D));
  generic_nmos I_2046(.D(I_2079_S), .G(I_2078_S), .S(VSS));
  generic_pmos I_2047(.D(I_2078_S), .G(I_1597_D), .S(VDD));
  generic_nmos I_2048(.D(I_2049_D), .G(I_2529_S), .S(I_2113_D));
  generic_pmos I_2049(.D(I_2049_D), .G(I_2305_S), .S(I_2113_D));
  generic_pmos I_205(.D(I_205_D), .G(I_205_G), .S(I_237_D));
  generic_nmos I_2050(.D(I_2050_D), .G(I_2050_G), .S(VSS));
  generic_pmos I_2051(.D(I_2051_D), .G(I_2147_S), .S(VDD));
  generic_nmos I_2052(.D(I_2053_D), .G(I_1831_S), .S(I_2053_S));
  generic_pmos I_2053(.D(I_2053_D), .G(I_1893_S), .S(I_2053_S));
  generic_nmos I_2054(.D(I_2055_D), .G(I_1893_S), .S(I_2055_S));
  generic_pmos I_2055(.D(I_2055_D), .G(I_1831_S), .S(I_2055_S));
  generic_nmos I_2056(.D(I_2056_D), .G(I_2056_G), .S(I_2056_S));
  generic_pmos I_2057(.D(I_2057_D), .G(I_2057_G), .S(I_2057_S));
  generic_nmos I_2058(.D(VSS), .G(I_2699_D), .S(I_2058_S));
  generic_pmos I_2059(.D(VDD), .G(I_2059_G), .S(I_2059_S));
  generic_nmos I_206(.D(I_206_D), .G(I_207_G), .S(I_238_D));
  generic_nmos I_2060(.D(I_2060_D), .G(I_2060_G), .S(I_2060_S));
  generic_pmos I_2061(.D(I_2061_D), .G(I_2061_G), .S(I_2061_S));
  generic_nmos I_2062(.D(I_2062_D), .G(I_2062_G), .S(VSS));
  generic_pmos I_2063(.D(I_2063_D), .G(I_2159_S), .S(VDD));
  generic_nmos I_2064(.D(I_2709_S), .G(I_2001_S), .S(I_2065_S));
  generic_pmos I_2065(.D(I_2709_S), .G(I_1969_D), .S(I_2065_S));
  generic_nmos I_2066(.D(I_2066_D), .G(I_2066_G), .S(I_2066_S));
  generic_pmos I_2067(.D(I_2067_D), .G(I_2067_G), .S(I_2067_S));
  generic_nmos I_2068(.D(I_2068_D), .G(I_2133_G), .S(VSS));
  generic_pmos I_2069(.D(I_2069_D), .G(I_1518_D), .S(VDD));
  generic_pmos I_207(.D(I_207_D), .G(I_207_G), .S(I_239_D));
  generic_nmos I_2070(.D(I_2071_D), .G(I_2103_D), .S(I_2071_S));
  generic_pmos I_2071(.D(I_2071_D), .G(I_2231_D), .S(I_2071_S));
  generic_nmos I_2072(.D(I_2073_D), .G(I_2007_D), .S(I_2169_D));
  generic_pmos I_2073(.D(I_2073_D), .G(I_1973_D), .S(I_2169_D));
  generic_nmos I_2074(.D(I_2074_D), .G(I_2071_D), .S(VSS));
  generic_pmos I_2075(.D(I_2075_D), .G(I_2171_S), .S(VDD));
  generic_nmos I_2076(.D(I_2076_D), .G(I_1917_D), .S(VSS));
  generic_pmos I_2077(.D(I_2077_D), .G(I_2013_D), .S(VDD));
  generic_nmos I_2078(.D(VSS), .G(I_1597_D), .S(I_2078_S));
  generic_pmos I_2079(.D(VDD), .G(I_2078_S), .S(I_2079_S));
  generic_nmos I_208(.D(I_208_D), .G(I_209_G), .S(I_240_D));
  generic_nmos I_2080(.D(I_2113_D), .G(I_2209_D), .S(I_2112_D));
  generic_pmos I_2081(.D(VDD), .G(I_2209_D), .S(I_2113_D));
  generic_nmos I_2082(.D(I_2115_D), .G(I_2083_G), .S(I_2114_D));
  generic_pmos I_2083(.D(VDD), .G(I_2083_G), .S(I_2115_D));
  generic_nmos I_2084(.D(I_2181_D), .G(I_2215_S), .S(VSS));
  generic_pmos I_2085(.D(I_2181_D), .G(I_2215_S), .S(VDD));
  generic_nmos I_2086(.D(I_2213_S), .G(I_2151_S), .S(I_2118_D));
  generic_pmos I_2087(.D(VDD), .G(I_2151_S), .S(I_2213_S));
  generic_nmos I_2088(.D(I_2088_D), .G(I_2089_G), .S(I_2120_D));
  generic_pmos I_2089(.D(I_2089_D), .G(I_2089_G), .S(I_2121_D));
  generic_pmos I_209(.D(I_209_D), .G(I_209_G), .S(I_241_D));
  generic_nmos I_2090(.D(I_2154_D), .G(I_2058_S), .S(VSS));
  generic_pmos I_2091(.D(I_2154_D), .G(I_2058_S), .S(I_2123_D));
  generic_nmos I_2092(.D(I_2092_D), .G(I_2093_G), .S(I_2124_D));
  generic_pmos I_2093(.D(I_2093_D), .G(I_2093_G), .S(I_2125_D));
  generic_nmos I_2094(.D(I_2127_D), .G(I_3271_S), .S(I_2126_D));
  generic_pmos I_2095(.D(VDD), .G(I_3271_S), .S(I_2127_D));
  generic_nmos I_2096(.D(I_2096_D), .G(I_2097_G), .S(I_2128_D));
  generic_pmos I_2097(.D(I_2097_D), .G(I_2097_G), .S(I_2129_D));
  generic_nmos I_2098(.D(I_2098_D), .G(I_2099_G), .S(I_2130_D));
  generic_pmos I_2099(.D(I_2099_D), .G(I_2099_G), .S(I_2131_D));
  generic_pmos I_21(.D(I_21_D), .G(I_21_G), .S(I_53_D));
  generic_nmos I_210(.D(I_210_D), .G(I_211_G), .S(I_242_D));
  generic_nmos I_2100(.D(VSS), .G(I_1518_D), .S(I_2132_D));
  generic_pmos I_2101(.D(I_2132_D), .G(I_1518_D), .S(I_2133_D));
  generic_nmos I_2102(.D(I_2103_D), .G(I_2231_D), .S(VSS));
  generic_pmos I_2103(.D(I_2103_D), .G(I_2231_D), .S(VDD));
  generic_nmos I_2104(.D(I_2105_D), .G(I_2073_D), .S(VSS));
  generic_pmos I_2105(.D(I_2105_D), .G(I_2073_D), .S(VDD));
  generic_nmos I_2106(.D(I_2139_D), .G(I_2169_D), .S(I_2138_D));
  generic_pmos I_2107(.D(VDD), .G(I_2169_D), .S(I_2139_D));
  generic_nmos I_2108(.D(I_2173_D), .G(I_2015_D), .S(I_2140_D));
  generic_pmos I_2109(.D(I_2173_D), .G(I_2015_D), .S(VDD));
  generic_pmos I_211(.D(I_211_D), .G(I_211_G), .S(I_243_D));
  generic_nmos I_2110(.D(I_2175_D), .G(I_3923_S), .S(I_2142_D));
  generic_pmos I_2111(.D(I_2175_D), .G(I_3923_S), .S(VDD));
  generic_nmos I_2112(.D(I_2112_D), .G(I_2113_G), .S(VSS));
  generic_pmos I_2113(.D(I_2113_D), .G(I_2113_G), .S(VDD));
  generic_nmos I_2114(.D(I_2114_D), .G(I_1033_D), .S(VSS));
  generic_pmos I_2115(.D(I_2115_D), .G(I_1033_D), .S(VDD));
  generic_nmos I_2116(.D(VSS), .G(I_1347_D), .S(I_2148_D));
  generic_pmos I_2117(.D(VDD), .G(I_1347_D), .S(I_2215_S));
  generic_nmos I_2118(.D(I_2118_D), .G(I_1347_D), .S(VSS));
  generic_pmos I_2119(.D(I_2213_S), .G(I_1347_D), .S(VDD));
  generic_nmos I_212(.D(VSS), .G(I_277_D), .S(I_245_D));
  generic_nmos I_2120(.D(I_2120_D), .G(I_2121_G), .S(I_2152_D));
  generic_pmos I_2121(.D(I_2121_D), .G(I_2121_G), .S(I_2153_D));
  generic_nmos I_2122(.D(VSS), .G(I_3562_D), .S(I_2154_D));
  generic_pmos I_2123(.D(I_2123_D), .G(I_3562_D), .S(I_2155_D));
  generic_nmos I_2124(.D(I_2124_D), .G(I_2125_G), .S(VSS));
  generic_pmos I_2125(.D(I_2125_D), .G(I_2125_G), .S(VDD));
  generic_nmos I_2126(.D(I_2126_D), .G(I_1997_D), .S(VSS));
  generic_pmos I_2127(.D(I_2127_D), .G(I_1997_D), .S(VDD));
  generic_nmos I_2128(.D(I_2128_D), .G(I_2129_G), .S(I_2160_D));
  generic_pmos I_2129(.D(I_2129_D), .G(I_2129_G), .S(I_2161_D));
  generic_pmos I_213(.D(VDD), .G(I_277_D), .S(I_245_D));
  generic_nmos I_2130(.D(I_2130_D), .G(I_2131_G), .S(I_2162_D));
  generic_pmos I_2131(.D(I_2131_D), .G(I_2131_G), .S(I_2163_D));
  generic_nmos I_2132(.D(I_2132_D), .G(I_2133_G), .S(VSS));
  generic_pmos I_2133(.D(I_2133_D), .G(I_2133_G), .S(VDD));
  generic_nmos I_2134(.D(VSS), .G(I_2135_G), .S(VSS));
  generic_pmos I_2135(.D(VDD), .G(I_2135_G), .S(VDD));
  generic_nmos I_2136(.D(VSS), .G(I_2105_D), .S(I_2169_D));
  generic_pmos I_2137(.D(VDD), .G(I_2105_D), .S(I_2169_D));
  generic_nmos I_2138(.D(I_2138_D), .G(I_1755_D), .S(VSS));
  generic_pmos I_2139(.D(I_2139_D), .G(I_1755_D), .S(VDD));
  generic_nmos I_214(.D(VSS), .G(I_311_D), .S(I_247_D));
  generic_nmos I_2140(.D(I_2140_D), .G(I_2175_D), .S(I_2172_D));
  generic_pmos I_2141(.D(VDD), .G(I_2175_D), .S(I_2173_D));
  generic_nmos I_2142(.D(I_2142_D), .G(I_2078_S), .S(I_2174_D));
  generic_pmos I_2143(.D(VDD), .G(I_2078_S), .S(I_2175_D));
  generic_nmos I_2144(.D(VSS), .G(I_2113_D), .S(I_2177_D));
  generic_pmos I_2145(.D(VDD), .G(I_2113_D), .S(I_2177_D));
  generic_nmos I_2146(.D(VSS), .G(I_1033_D), .S(I_2147_S));
  generic_pmos I_2147(.D(VDD), .G(I_1033_D), .S(I_2147_S));
  generic_nmos I_2148(.D(I_2148_D), .G(I_2213_D), .S(I_2215_S));
  generic_pmos I_2149(.D(I_2215_S), .G(I_2213_D), .S(VDD));
  generic_pmos I_215(.D(VDD), .G(I_311_D), .S(I_247_D));
  generic_nmos I_2150(.D(VSS), .G(I_2215_D), .S(I_2151_S));
  generic_pmos I_2151(.D(VDD), .G(I_2215_D), .S(I_2151_S));
  generic_nmos I_2152(.D(I_2152_D), .G(I_2153_G), .S(I_2152_S));
  generic_pmos I_2153(.D(I_2153_D), .G(I_2153_G), .S(I_2153_S));
  generic_nmos I_2154(.D(I_2154_D), .G(I_2539_S), .S(VSS));
  generic_pmos I_2155(.D(I_2155_D), .G(I_2539_S), .S(VDD));
  generic_nmos I_2156(.D(VSS), .G(I_873_D), .S(I_2157_S));
  generic_pmos I_2157(.D(VDD), .G(I_873_D), .S(I_2157_S));
  generic_nmos I_2158(.D(VSS), .G(I_1997_D), .S(I_2159_S));
  generic_pmos I_2159(.D(VDD), .G(I_1997_D), .S(I_2159_S));
  generic_nmos I_216(.D(VSS), .G(I_153_D), .S(I_281_D));
  generic_nmos I_2160(.D(I_2160_D), .G(I_2161_G), .S(I_2160_S));
  generic_pmos I_2161(.D(I_2161_D), .G(I_2161_G), .S(I_2161_S));
  generic_nmos I_2162(.D(I_2162_D), .G(I_2163_G), .S(I_2162_S));
  generic_pmos I_2163(.D(I_2163_D), .G(I_2163_G), .S(I_2163_S));
  generic_nmos I_2164(.D(VSS), .G(I_2132_D), .S(I_2165_S));
  generic_pmos I_2165(.D(VDD), .G(I_2132_D), .S(I_2165_S));
  generic_nmos I_2166(.D(VSS), .G(I_2071_S), .S(I_2167_S));
  generic_pmos I_2167(.D(VDD), .G(I_2071_S), .S(I_2167_S));
  generic_nmos I_2168(.D(I_2169_D), .G(I_2105_D), .S(VSS));
  generic_pmos I_2169(.D(I_2169_D), .G(I_2105_D), .S(VDD));
  generic_pmos I_217(.D(VDD), .G(I_153_D), .S(I_281_D));
  generic_nmos I_2170(.D(VSS), .G(I_1755_D), .S(I_2171_S));
  generic_pmos I_2171(.D(VDD), .G(I_1755_D), .S(I_2171_S));
  generic_nmos I_2172(.D(I_2172_D), .G(I_2335_D), .S(VSS));
  generic_pmos I_2173(.D(I_2173_D), .G(I_2335_D), .S(VDD));
  generic_nmos I_2174(.D(I_2174_D), .G(I_2239_S), .S(VSS));
  generic_pmos I_2175(.D(I_2175_D), .G(I_2239_S), .S(VDD));
  generic_nmos I_2176(.D(I_2177_D), .G(I_2529_S), .S(I_2209_D));
  generic_pmos I_2177(.D(I_2177_D), .G(I_2305_S), .S(I_2209_D));
  generic_nmos I_2178(.D(I_2211_D), .G(I_2213_S), .S(I_2210_D));
  generic_pmos I_2179(.D(VDD), .G(I_2053_S), .S(I_2211_D));
  generic_nmos I_218(.D(I_251_S), .G(I_347_D), .S(VSS));
  generic_nmos I_2180(.D(I_2181_D), .G(I_2053_S), .S(I_2213_D));
  generic_pmos I_2181(.D(I_2181_D), .G(I_1991_S), .S(I_2213_D));
  generic_nmos I_2182(.D(I_2213_S), .G(I_1991_S), .S(I_2215_D));
  generic_pmos I_2183(.D(I_2213_S), .G(I_2053_S), .S(I_2215_D));
  generic_nmos I_2184(.D(I_2184_D), .G(I_2184_G), .S(I_2216_D));
  generic_pmos I_2185(.D(I_2185_D), .G(I_2216_G), .S(I_2217_D));
  generic_nmos I_2186(.D(I_2219_S), .G(I_2154_D), .S(VSS));
  generic_pmos I_2187(.D(I_2187_D), .G(I_2218_G), .S(VDD));
  generic_nmos I_2188(.D(VSS), .G(I_2317_S), .S(I_2253_D));
  generic_pmos I_2189(.D(VDD), .G(I_2317_S), .S(I_2253_D));
  generic_pmos I_219(.D(I_251_S), .G(I_347_D), .S(VDD));
  generic_nmos I_2190(.D(I_2190_D), .G(I_2190_G), .S(I_2222_D));
  generic_pmos I_2191(.D(I_2191_D), .G(I_2222_G), .S(I_2223_D));
  generic_nmos I_2192(.D(I_2225_D), .G(I_1999_D), .S(I_2224_D));
  generic_pmos I_2193(.D(VDD), .G(I_2319_D), .S(I_2225_D));
  generic_nmos I_2194(.D(I_2194_D), .G(I_2194_G), .S(I_2226_D));
  generic_pmos I_2195(.D(I_2195_D), .G(I_2226_G), .S(I_2227_D));
  generic_nmos I_2196(.D(VSS), .G(I_2132_D), .S(I_2711_S));
  generic_pmos I_2197(.D(I_2197_D), .G(I_2228_G), .S(I_2711_S));
  generic_nmos I_2198(.D(I_2231_D), .G(I_2071_S), .S(I_2231_S));
  generic_pmos I_2199(.D(I_2199_D), .G(I_2167_S), .S(I_2231_D));
  generic_nmos I_22(.D(I_2521_D), .G(I_23_G), .S(VSS));
  generic_nmos I_220(.D(I_220_D), .G(I_159_S), .S(VSS));
  generic_nmos I_2200(.D(I_2201_D), .G(I_1973_D), .S(I_2233_D));
  generic_pmos I_2201(.D(I_2201_D), .G(I_2007_D), .S(I_2233_D));
  generic_nmos I_2202(.D(VSS), .G(I_2267_D), .S(I_2234_D));
  generic_pmos I_2203(.D(VDD), .G(I_2549_D), .S(I_2235_D));
  generic_nmos I_2204(.D(VSS), .G(I_2269_D), .S(I_2236_D));
  generic_pmos I_2205(.D(VDD), .G(I_2173_D), .S(I_2237_D));
  generic_nmos I_2206(.D(I_2239_S), .G(I_2238_S), .S(VSS));
  generic_pmos I_2207(.D(I_2238_S), .G(I_1821_D), .S(VDD));
  generic_nmos I_2208(.D(I_2209_D), .G(I_2305_S), .S(I_2209_S));
  generic_pmos I_2209(.D(I_2209_D), .G(I_2529_S), .S(I_2209_S));
  generic_pmos I_221(.D(I_285_D), .G(I_159_S), .S(VDD));
  generic_nmos I_2210(.D(I_2210_D), .G(I_2053_S), .S(VSS));
  generic_pmos I_2211(.D(I_2211_D), .G(I_2213_S), .S(VDD));
  generic_nmos I_2212(.D(I_2213_D), .G(I_1991_S), .S(I_2213_S));
  generic_pmos I_2213(.D(I_2213_D), .G(I_2053_S), .S(I_2213_S));
  generic_nmos I_2214(.D(I_2215_D), .G(I_2053_S), .S(I_2215_S));
  generic_pmos I_2215(.D(I_2215_D), .G(I_1991_S), .S(I_2215_S));
  generic_nmos I_2216(.D(I_2216_D), .G(I_2216_G), .S(I_2216_S));
  generic_pmos I_2217(.D(I_2217_D), .G(I_2217_G), .S(I_2217_S));
  generic_nmos I_2218(.D(VSS), .G(I_2218_G), .S(I_2218_S));
  generic_pmos I_2219(.D(VDD), .G(I_2154_D), .S(I_2219_S));
  generic_nmos I_222(.D(I_222_D), .G(I_223_G), .S(I_254_D));
  generic_nmos I_2220(.D(I_2253_D), .G(I_2317_S), .S(VSS));
  generic_pmos I_2221(.D(I_2253_D), .G(I_2317_S), .S(VDD));
  generic_nmos I_2222(.D(I_2222_D), .G(I_2222_G), .S(I_2222_S));
  generic_pmos I_2223(.D(I_2223_D), .G(I_2223_G), .S(I_2223_S));
  generic_nmos I_2224(.D(I_2224_D), .G(I_2319_D), .S(VSS));
  generic_pmos I_2225(.D(I_2225_D), .G(I_1999_D), .S(VDD));
  generic_nmos I_2226(.D(I_2226_D), .G(I_2226_G), .S(I_2226_S));
  generic_pmos I_2227(.D(I_2227_D), .G(I_2227_G), .S(I_2227_S));
  generic_nmos I_2228(.D(I_2711_S), .G(I_2228_G), .S(I_2228_S));
  generic_pmos I_2229(.D(I_2711_S), .G(I_2069_D), .S(VDD));
  generic_pmos I_223(.D(I_223_D), .G(I_223_G), .S(I_255_D));
  generic_nmos I_2230(.D(I_2231_S), .G(I_2167_S), .S(VSS));
  generic_pmos I_2231(.D(I_2231_D), .G(I_2167_S), .S(I_2231_S));
  generic_nmos I_2232(.D(I_2233_D), .G(I_2007_D), .S(I_2329_D));
  generic_pmos I_2233(.D(I_2233_D), .G(I_1973_D), .S(I_2329_D));
  generic_nmos I_2234(.D(I_2234_D), .G(I_2549_D), .S(I_2235_D));
  generic_pmos I_2235(.D(I_2235_D), .G(I_2267_D), .S(VDD));
  generic_nmos I_2236(.D(I_2236_D), .G(I_2173_D), .S(I_2237_D));
  generic_pmos I_2237(.D(I_2237_D), .G(I_2269_D), .S(VDD));
  generic_nmos I_2238(.D(VSS), .G(I_1821_D), .S(I_2238_S));
  generic_pmos I_2239(.D(VDD), .G(I_2238_S), .S(I_2239_S));
  generic_nmos I_224(.D(I_224_D), .G(I_289_D), .S(VSS));
  generic_nmos I_2240(.D(I_2529_S), .G(I_2241_G), .S(I_2272_D));
  generic_pmos I_2241(.D(VDD), .G(I_2241_G), .S(I_2529_S));
  generic_nmos I_2242(.D(I_2275_D), .G(I_2311_S), .S(I_2274_D));
  generic_pmos I_2243(.D(VDD), .G(I_2311_S), .S(I_2275_D));
  generic_nmos I_2244(.D(I_2341_D), .G(I_2375_S), .S(VSS));
  generic_pmos I_2245(.D(I_2341_D), .G(I_2375_S), .S(VDD));
  generic_nmos I_2246(.D(I_2373_S), .G(I_2311_S), .S(I_2278_D));
  generic_pmos I_2247(.D(VDD), .G(I_2311_S), .S(I_2373_S));
  generic_nmos I_2248(.D(I_2248_D), .G(I_2249_G), .S(I_2280_D));
  generic_pmos I_2249(.D(I_2249_D), .G(I_2249_G), .S(I_2281_D));
  generic_pmos I_225(.D(I_225_D), .G(I_289_D), .S(VDD));
  generic_nmos I_2250(.D(I_3499_D), .G(I_873_D), .S(I_2282_D));
  generic_pmos I_2251(.D(VDD), .G(I_873_D), .S(I_3499_D));
  generic_nmos I_2252(.D(I_2253_D), .G(I_2317_S), .S(VSS));
  generic_pmos I_2253(.D(I_2253_D), .G(I_2317_S), .S(VDD));
  generic_nmos I_2254(.D(I_2254_D), .G(I_2255_G), .S(VSS));
  generic_pmos I_2255(.D(I_2255_D), .G(I_2255_G), .S(VDD));
  generic_nmos I_2256(.D(VSS), .G(I_1999_D), .S(I_2288_D));
  generic_pmos I_2257(.D(I_2288_D), .G(I_1999_D), .S(I_2289_D));
  generic_nmos I_2258(.D(I_2258_D), .G(I_2259_G), .S(I_2290_D));
  generic_pmos I_2259(.D(I_2259_D), .G(I_2259_G), .S(I_2291_D));
  generic_nmos I_226(.D(I_226_D), .G(I_355_D), .S(I_227_D));
  generic_nmos I_2260(.D(I_2549_S), .G(I_2165_S), .S(I_2292_D));
  generic_pmos I_2261(.D(VDD), .G(I_2165_S), .S(I_2549_S));
  generic_nmos I_2262(.D(I_2263_D), .G(I_2231_S), .S(VSS));
  generic_pmos I_2263(.D(I_2263_D), .G(I_2231_S), .S(VDD));
  generic_nmos I_2264(.D(I_2265_D), .G(I_2233_D), .S(VSS));
  generic_pmos I_2265(.D(I_2265_D), .G(I_2233_D), .S(VDD));
  generic_nmos I_2266(.D(I_2267_D), .G(I_1755_D), .S(VSS));
  generic_pmos I_2267(.D(I_2267_D), .G(I_1755_D), .S(VDD));
  generic_nmos I_2268(.D(I_2269_D), .G(I_2009_D), .S(VSS));
  generic_pmos I_2269(.D(I_2269_D), .G(I_2009_D), .S(VDD));
  generic_pmos I_227(.D(I_227_D), .G(I_355_D), .S(VDD));
  generic_nmos I_2270(.D(I_2335_D), .G(I_2079_S), .S(I_2302_D));
  generic_pmos I_2271(.D(I_2335_D), .G(I_2079_S), .S(VDD));
  generic_nmos I_2272(.D(I_2272_D), .G(I_2305_S), .S(VSS));
  generic_pmos I_2273(.D(I_2529_S), .G(I_2305_S), .S(VDD));
  generic_nmos I_2274(.D(I_2274_D), .G(I_2211_D), .S(VSS));
  generic_pmos I_2275(.D(I_2275_D), .G(I_2211_D), .S(VDD));
  generic_nmos I_2276(.D(VSS), .G(I_1347_D), .S(I_2308_D));
  generic_pmos I_2277(.D(VDD), .G(I_1347_D), .S(I_2375_S));
  generic_nmos I_2278(.D(I_2278_D), .G(I_1347_D), .S(VSS));
  generic_pmos I_2279(.D(I_2373_S), .G(I_1347_D), .S(VDD));
  generic_nmos I_228(.D(VSS), .G(I_293_D), .S(I_229_S));
  generic_nmos I_2280(.D(I_2280_D), .G(I_2281_G), .S(I_2312_D));
  generic_pmos I_2281(.D(I_2281_D), .G(I_2281_G), .S(I_2313_D));
  generic_nmos I_2282(.D(I_2282_D), .G(I_2219_S), .S(VSS));
  generic_pmos I_2283(.D(I_3499_D), .G(I_2219_S), .S(VDD));
  generic_nmos I_2284(.D(VSS), .G(I_2285_G), .S(VSS));
  generic_pmos I_2285(.D(VDD), .G(I_2285_G), .S(VDD));
  generic_nmos I_2286(.D(VSS), .G(I_2383_D), .S(I_2318_D));
  generic_pmos I_2287(.D(VDD), .G(I_2383_D), .S(I_2319_D));
  generic_nmos I_2288(.D(I_2288_D), .G(I_2319_D), .S(VSS));
  generic_pmos I_2289(.D(I_2289_D), .G(I_2319_D), .S(VDD));
  generic_pmos I_229(.D(VDD), .G(I_293_D), .S(I_229_S));
  generic_nmos I_2290(.D(I_2290_D), .G(I_2291_G), .S(I_2322_D));
  generic_pmos I_2291(.D(I_2291_D), .G(I_2291_G), .S(I_2323_D));
  generic_nmos I_2292(.D(I_2292_D), .G(I_2069_D), .S(VSS));
  generic_pmos I_2293(.D(I_2549_S), .G(I_2069_D), .S(VDD));
  generic_nmos I_2294(.D(VSS), .G(I_2295_G), .S(VSS));
  generic_pmos I_2295(.D(VDD), .G(I_2295_G), .S(VDD));
  generic_nmos I_2296(.D(VSS), .G(I_2265_D), .S(I_2329_D));
  generic_pmos I_2297(.D(VDD), .G(I_2265_D), .S(I_2329_D));
  generic_nmos I_2298(.D(VSS), .G(I_1755_D), .S(I_2330_D));
  generic_pmos I_2299(.D(VDD), .G(I_1755_D), .S(I_2331_D));
  generic_pmos I_23(.D(I_2521_D), .G(I_23_G), .S(VDD));
  generic_nmos I_230(.D(I_230_D), .G(I_295_D), .S(I_293_S));
  generic_nmos I_2300(.D(VSS), .G(I_2009_D), .S(I_2332_D));
  generic_pmos I_2301(.D(VDD), .G(I_2009_D), .S(I_2333_D));
  generic_nmos I_2302(.D(I_2302_D), .G(I_2238_S), .S(I_2334_D));
  generic_pmos I_2303(.D(VDD), .G(I_2238_S), .S(I_2335_D));
  generic_nmos I_2304(.D(VSS), .G(I_2369_D), .S(I_2305_S));
  generic_pmos I_2305(.D(VDD), .G(I_2369_D), .S(I_2305_S));
  generic_nmos I_2306(.D(VSS), .G(I_2307_G), .S(I_2306_S));
  generic_pmos I_2307(.D(VDD), .G(I_2307_G), .S(I_2307_S));
  generic_nmos I_2308(.D(I_2308_D), .G(I_2373_D), .S(I_2375_S));
  generic_pmos I_2309(.D(I_2375_S), .G(I_2373_D), .S(VDD));
  generic_pmos I_231(.D(I_293_S), .G(I_295_D), .S(VDD));
  generic_nmos I_2310(.D(VSS), .G(I_2375_D), .S(I_2311_S));
  generic_pmos I_2311(.D(VDD), .G(I_2375_D), .S(I_2311_S));
  generic_nmos I_2312(.D(I_2312_D), .G(I_2313_G), .S(I_2312_S));
  generic_pmos I_2313(.D(I_2313_D), .G(I_2313_G), .S(I_2313_S));
  generic_nmos I_2314(.D(VSS), .G(I_2315_G), .S(I_2314_S));
  generic_pmos I_2315(.D(VDD), .G(I_2315_G), .S(I_2315_S));
  generic_nmos I_2316(.D(VSS), .G(I_3499_D), .S(I_2317_S));
  generic_pmos I_2317(.D(VDD), .G(I_3499_D), .S(I_2317_S));
  generic_nmos I_2318(.D(I_2318_D), .G(I_2447_D), .S(I_2319_D));
  generic_pmos I_2319(.D(I_2319_D), .G(I_2447_D), .S(VDD));
  generic_nmos I_232(.D(I_232_D), .G(I_233_G), .S(I_232_S));
  generic_nmos I_2320(.D(VSS), .G(I_2288_D), .S(I_2321_S));
  generic_pmos I_2321(.D(VDD), .G(I_2288_D), .S(I_2321_S));
  generic_nmos I_2322(.D(I_2322_D), .G(I_2323_G), .S(I_2322_S));
  generic_pmos I_2323(.D(I_2323_D), .G(I_2323_G), .S(I_2323_S));
  generic_nmos I_2324(.D(VSS), .G(I_2549_S), .S(I_2517_D));
  generic_pmos I_2325(.D(VDD), .G(I_2549_S), .S(I_2517_D));
  generic_nmos I_2326(.D(VSS), .G(I_2263_D), .S(I_2389_S));
  generic_pmos I_2327(.D(VDD), .G(I_2263_D), .S(I_2389_S));
  generic_nmos I_2328(.D(I_2329_D), .G(I_2265_D), .S(VSS));
  generic_pmos I_2329(.D(I_2329_D), .G(I_2265_D), .S(VDD));
  generic_pmos I_233(.D(I_233_D), .G(I_233_G), .S(I_233_S));
  generic_nmos I_2330(.D(I_2330_D), .G(I_2329_D), .S(I_2331_D));
  generic_pmos I_2331(.D(I_2331_D), .G(I_2329_D), .S(VDD));
  generic_nmos I_2332(.D(I_2332_D), .G(I_2395_D), .S(I_2333_D));
  generic_pmos I_2333(.D(I_2333_D), .G(I_2395_D), .S(VDD));
  generic_nmos I_2334(.D(I_2334_D), .G(VDD), .S(VSS));
  generic_pmos I_2335(.D(I_2335_D), .G(VDD), .S(VDD));
  generic_nmos I_2336(.D(I_2529_S), .G(I_2625_S), .S(I_2369_D));
  generic_pmos I_2337(.D(I_2529_S), .G(I_2657_D), .S(I_2369_D));
  generic_nmos I_2338(.D(VSS), .G(I_2632_D), .S(I_2371_S));
  generic_pmos I_2339(.D(VDD), .G(I_2370_G), .S(I_2371_D));
  generic_nmos I_234(.D(I_234_D), .G(I_618_S), .S(VSS));
  generic_nmos I_2340(.D(I_2341_D), .G(I_2213_S), .S(I_2373_D));
  generic_pmos I_2341(.D(I_2341_D), .G(I_2151_S), .S(I_2373_D));
  generic_nmos I_2342(.D(I_2373_S), .G(I_2151_S), .S(I_2375_D));
  generic_pmos I_2343(.D(I_2373_S), .G(I_2213_S), .S(I_2375_D));
  generic_nmos I_2344(.D(I_2344_D), .G(I_2344_G), .S(I_2376_D));
  generic_pmos I_2345(.D(I_2345_D), .G(I_2376_G), .S(I_2377_D));
  generic_nmos I_2346(.D(VSS), .G(I_3499_D), .S(I_2379_S));
  generic_pmos I_2347(.D(VDD), .G(I_3337_D), .S(I_2379_D));
  generic_nmos I_2348(.D(I_2348_D), .G(I_2348_G), .S(VSS));
  generic_pmos I_2349(.D(VDD), .G(I_3337_D), .S(VDD));
  generic_pmos I_235(.D(I_235_D), .G(I_618_S), .S(VDD));
  generic_nmos I_2350(.D(I_2383_D), .G(I_2479_S), .S(I_2382_D));
  generic_pmos I_2351(.D(VDD), .G(I_3111_S), .S(I_2383_D));
  generic_nmos I_2352(.D(VSS), .G(I_2288_D), .S(I_3185_S));
  generic_pmos I_2353(.D(I_2353_D), .G(I_2384_G), .S(I_3185_S));
  generic_nmos I_2354(.D(I_2354_D), .G(I_2354_G), .S(I_2386_D));
  generic_pmos I_2355(.D(I_2355_D), .G(I_2386_G), .S(I_2387_D));
  generic_nmos I_2356(.D(I_2711_S), .G(I_2517_D), .S(I_2389_S));
  generic_pmos I_2357(.D(I_2357_D), .G(I_2388_G), .S(I_2711_S));
  generic_nmos I_2358(.D(I_2391_D), .G(I_1265_D), .S(I_2390_D));
  generic_pmos I_2359(.D(VDD), .G(I_2311_S), .S(I_2391_D));
  generic_nmos I_236(.D(I_236_D), .G(I_237_G), .S(I_236_S));
  generic_nmos I_2360(.D(I_2361_D), .G(I_1973_D), .S(I_2393_D));
  generic_pmos I_2361(.D(I_2361_D), .G(I_2007_D), .S(I_2393_D));
  generic_nmos I_2362(.D(I_2395_D), .G(I_2331_D), .S(I_2394_D));
  generic_pmos I_2363(.D(VDD), .G(I_2235_D), .S(I_2395_D));
  generic_nmos I_2364(.D(I_2397_D), .G(I_2333_D), .S(I_2396_D));
  generic_pmos I_2365(.D(VDD), .G(I_2237_D), .S(I_2397_D));
  generic_nmos I_2366(.D(VSS), .G(I_2397_D), .S(I_2399_D));
  generic_pmos I_2367(.D(VDD), .G(I_2397_D), .S(I_2399_D));
  generic_nmos I_2368(.D(I_2369_D), .G(I_2657_D), .S(I_2433_D));
  generic_pmos I_2369(.D(I_2369_D), .G(I_2625_S), .S(I_2433_D));
  generic_pmos I_237(.D(I_237_D), .G(I_237_G), .S(I_237_S));
  generic_nmos I_2370(.D(I_2371_S), .G(I_2370_G), .S(VSS));
  generic_pmos I_2371(.D(I_2371_D), .G(I_2632_D), .S(I_2371_S));
  generic_nmos I_2372(.D(I_2373_D), .G(I_2151_S), .S(I_2373_S));
  generic_pmos I_2373(.D(I_2373_D), .G(I_2213_S), .S(I_2373_S));
  generic_nmos I_2374(.D(I_2375_D), .G(I_2213_S), .S(I_2375_S));
  generic_pmos I_2375(.D(I_2375_D), .G(I_2151_S), .S(I_2375_S));
  generic_nmos I_2376(.D(I_2376_D), .G(I_2376_G), .S(I_2376_S));
  generic_pmos I_2377(.D(I_2377_D), .G(I_2377_G), .S(I_2377_S));
  generic_nmos I_2378(.D(I_2379_S), .G(I_3337_D), .S(VSS));
  generic_pmos I_2379(.D(I_2379_D), .G(I_3499_D), .S(I_2379_S));
  generic_nmos I_238(.D(I_238_D), .G(I_239_G), .S(I_238_S));
  generic_nmos I_2380(.D(VSS), .G(I_3337_D), .S(VSS));
  generic_pmos I_2381(.D(VDD), .G(I_2381_G), .S(I_2381_S));
  generic_nmos I_2382(.D(I_2382_D), .G(I_3111_S), .S(VSS));
  generic_pmos I_2383(.D(I_2383_D), .G(I_2479_S), .S(VDD));
  generic_nmos I_2384(.D(I_3185_S), .G(I_2384_G), .S(I_2384_S));
  generic_pmos I_2385(.D(I_3185_S), .G(I_2225_D), .S(VDD));
  generic_nmos I_2386(.D(I_2386_D), .G(I_2386_G), .S(I_2386_S));
  generic_pmos I_2387(.D(I_2387_D), .G(I_2387_G), .S(I_2387_S));
  generic_nmos I_2388(.D(I_2389_S), .G(I_2388_G), .S(I_2388_S));
  generic_pmos I_2389(.D(I_2711_S), .G(I_2549_S), .S(I_2389_S));
  generic_pmos I_239(.D(I_239_D), .G(I_239_G), .S(I_239_S));
  generic_nmos I_2390(.D(I_2390_D), .G(I_2311_S), .S(VSS));
  generic_pmos I_2391(.D(I_2391_D), .G(I_1265_D), .S(VDD));
  generic_nmos I_2392(.D(I_2393_D), .G(I_2007_D), .S(I_2489_D));
  generic_pmos I_2393(.D(I_2393_D), .G(I_1973_D), .S(I_2489_D));
  generic_nmos I_2394(.D(I_2394_D), .G(I_2235_D), .S(VSS));
  generic_pmos I_2395(.D(I_2395_D), .G(I_2331_D), .S(VDD));
  generic_nmos I_2396(.D(I_2396_D), .G(I_2237_D), .S(VSS));
  generic_pmos I_2397(.D(I_2397_D), .G(I_2333_D), .S(VDD));
  generic_nmos I_2398(.D(I_2399_D), .G(I_2397_D), .S(VSS));
  generic_pmos I_2399(.D(I_2399_D), .G(I_2397_D), .S(VDD));
  generic_nmos I_24(.D(I_24_D), .G(I_25_G), .S(I_56_D));
  generic_nmos I_240(.D(I_240_D), .G(I_241_G), .S(I_240_S));
  generic_nmos I_2400(.D(I_2433_D), .G(I_2529_D), .S(I_2432_D));
  generic_pmos I_2401(.D(VDD), .G(I_2529_D), .S(I_2433_D));
  generic_nmos I_2402(.D(I_2402_D), .G(I_2403_G), .S(I_2434_D));
  generic_pmos I_2403(.D(I_2403_D), .G(I_2403_G), .S(I_2435_D));
  generic_nmos I_2404(.D(I_2501_D), .G(I_2535_S), .S(VSS));
  generic_pmos I_2405(.D(I_2501_D), .G(I_2535_S), .S(VDD));
  generic_nmos I_2406(.D(I_2533_S), .G(I_2471_S), .S(I_2438_D));
  generic_pmos I_2407(.D(VDD), .G(I_2471_S), .S(I_2533_S));
  generic_nmos I_2408(.D(I_2408_D), .G(I_2409_G), .S(I_2440_D));
  generic_pmos I_2409(.D(I_2409_D), .G(I_2409_G), .S(I_2441_D));
  generic_pmos I_241(.D(I_241_D), .G(I_241_G), .S(I_241_S));
  generic_nmos I_2410(.D(I_2410_D), .G(I_2411_G), .S(I_2442_D));
  generic_pmos I_2411(.D(I_2411_D), .G(I_2411_G), .S(I_2443_D));
  generic_nmos I_2412(.D(I_2412_D), .G(I_2413_G), .S(I_2444_D));
  generic_pmos I_2413(.D(I_2413_D), .G(I_2413_G), .S(I_2445_D));
  generic_nmos I_2414(.D(I_2447_D), .G(I_3337_D), .S(I_2446_D));
  generic_pmos I_2415(.D(VDD), .G(I_3337_D), .S(I_2447_D));
  generic_nmos I_2416(.D(I_2705_S), .G(I_2321_S), .S(I_2448_D));
  generic_pmos I_2417(.D(VDD), .G(I_2321_S), .S(I_2705_S));
  generic_nmos I_2418(.D(I_2418_D), .G(I_2419_G), .S(I_2450_D));
  generic_pmos I_2419(.D(I_2419_D), .G(I_2419_G), .S(I_2451_D));
  generic_nmos I_242(.D(I_242_D), .G(I_243_G), .S(I_242_S));
  generic_nmos I_2420(.D(I_2420_D), .G(I_2421_G), .S(I_2453_D));
  generic_pmos I_2421(.D(I_2421_D), .G(I_2421_G), .S(I_2453_D));
  generic_nmos I_2422(.D(VSS), .G(I_1265_D), .S(I_2454_D));
  generic_pmos I_2423(.D(I_2454_D), .G(I_1265_D), .S(I_2455_D));
  generic_nmos I_2424(.D(I_2425_D), .G(I_2393_D), .S(VSS));
  generic_pmos I_2425(.D(I_2425_D), .G(I_2393_D), .S(VDD));
  generic_nmos I_2426(.D(I_2427_D), .G(I_1755_D), .S(VSS));
  generic_pmos I_2427(.D(I_2427_D), .G(I_1755_D), .S(VDD));
  generic_nmos I_2428(.D(I_2429_D), .G(I_2009_D), .S(VSS));
  generic_pmos I_2429(.D(I_2429_D), .G(I_2009_D), .S(VDD));
  generic_pmos I_243(.D(I_243_D), .G(I_243_G), .S(I_243_S));
  generic_nmos I_2430(.D(I_2495_D), .G(I_3036_S), .S(I_2462_D));
  generic_pmos I_2431(.D(I_2495_D), .G(I_3036_S), .S(VDD));
  generic_nmos I_2432(.D(I_2432_D), .G(I_2433_G), .S(VSS));
  generic_pmos I_2433(.D(I_2433_D), .G(I_2433_G), .S(VDD));
  generic_nmos I_2434(.D(I_2434_D), .G(I_2435_G), .S(I_2466_D));
  generic_pmos I_2435(.D(I_2435_D), .G(I_2435_G), .S(I_2467_D));
  generic_nmos I_2436(.D(VSS), .G(I_3241_D), .S(I_2468_D));
  generic_pmos I_2437(.D(VDD), .G(I_3241_D), .S(I_2535_S));
  generic_nmos I_2438(.D(I_2438_D), .G(I_3241_D), .S(VSS));
  generic_pmos I_2439(.D(I_2533_S), .G(I_3241_D), .S(VDD));
  generic_nmos I_244(.D(I_245_D), .G(I_277_D), .S(VSS));
  generic_nmos I_2440(.D(I_2440_D), .G(I_2441_G), .S(I_2472_D));
  generic_pmos I_2441(.D(I_2441_D), .G(I_2441_G), .S(I_2473_D));
  generic_nmos I_2442(.D(I_2442_D), .G(I_2443_G), .S(I_2474_D));
  generic_pmos I_2443(.D(I_2443_D), .G(I_2443_G), .S(I_2475_D));
  generic_nmos I_2444(.D(I_2444_D), .G(I_2445_G), .S(I_2476_D));
  generic_pmos I_2445(.D(I_2445_D), .G(I_2445_G), .S(I_2477_D));
  generic_nmos I_2446(.D(I_2446_D), .G(I_2253_D), .S(VSS));
  generic_pmos I_2447(.D(I_2447_D), .G(I_2253_D), .S(VDD));
  generic_nmos I_2448(.D(I_2448_D), .G(I_2225_D), .S(VSS));
  generic_pmos I_2449(.D(I_2705_S), .G(I_2225_D), .S(VDD));
  generic_pmos I_245(.D(I_245_D), .G(I_277_D), .S(VDD));
  generic_nmos I_2450(.D(I_2450_D), .G(I_2451_G), .S(I_2482_D));
  generic_pmos I_2451(.D(I_2451_D), .G(I_2451_G), .S(I_2483_D));
  generic_nmos I_2452(.D(I_2453_D), .G(I_2389_S), .S(VSS));
  generic_pmos I_2453(.D(I_2453_D), .G(I_2389_S), .S(VDD));
  generic_nmos I_2454(.D(I_2454_D), .G(I_2311_S), .S(VSS));
  generic_pmos I_2455(.D(I_2455_D), .G(I_2311_S), .S(VDD));
  generic_nmos I_2456(.D(VSS), .G(I_2425_D), .S(I_2489_D));
  generic_pmos I_2457(.D(VDD), .G(I_2425_D), .S(I_2489_D));
  generic_nmos I_2458(.D(VSS), .G(I_1755_D), .S(I_2490_D));
  generic_pmos I_2459(.D(VDD), .G(I_1755_D), .S(I_2491_D));
  generic_nmos I_246(.D(I_247_D), .G(I_311_D), .S(VSS));
  generic_nmos I_2460(.D(VSS), .G(I_2009_D), .S(I_2492_D));
  generic_pmos I_2461(.D(VDD), .G(I_2009_D), .S(I_2493_D));
  generic_nmos I_2462(.D(I_2462_D), .G(I_2718_S), .S(I_2494_D));
  generic_pmos I_2463(.D(VDD), .G(I_2718_S), .S(I_2495_D));
  generic_nmos I_2464(.D(VSS), .G(I_2433_D), .S(I_2497_D));
  generic_pmos I_2465(.D(VDD), .G(I_2433_D), .S(I_2497_D));
  generic_nmos I_2466(.D(I_2466_D), .G(I_2467_G), .S(I_2466_S));
  generic_pmos I_2467(.D(I_2467_D), .G(I_2467_G), .S(I_2467_S));
  generic_nmos I_2468(.D(I_2468_D), .G(I_2533_D), .S(I_2535_S));
  generic_pmos I_2469(.D(I_2535_S), .G(I_2533_D), .S(VDD));
  generic_pmos I_247(.D(I_247_D), .G(I_311_D), .S(VDD));
  generic_nmos I_2470(.D(VSS), .G(I_2535_D), .S(I_2471_S));
  generic_pmos I_2471(.D(VDD), .G(I_2535_D), .S(I_2471_S));
  generic_nmos I_2472(.D(I_2472_D), .G(I_2473_G), .S(I_2472_S));
  generic_pmos I_2473(.D(I_2473_D), .G(I_2473_G), .S(I_2473_S));
  generic_nmos I_2474(.D(I_2474_D), .G(I_2475_G), .S(I_2474_S));
  generic_pmos I_2475(.D(I_2475_D), .G(I_2475_G), .S(I_2475_S));
  generic_nmos I_2476(.D(I_2476_D), .G(I_2477_G), .S(I_2476_S));
  generic_pmos I_2477(.D(I_2477_D), .G(I_2477_G), .S(I_2477_S));
  generic_nmos I_2478(.D(VSS), .G(I_2253_D), .S(I_2479_S));
  generic_pmos I_2479(.D(VDD), .G(I_2253_D), .S(I_2479_S));
  generic_nmos I_248(.D(I_281_D), .G(I_153_D), .S(VSS));
  generic_nmos I_2480(.D(VSS), .G(I_2705_S), .S(I_2673_D));
  generic_pmos I_2481(.D(VDD), .G(I_2705_S), .S(I_2673_D));
  generic_nmos I_2482(.D(I_2482_D), .G(I_2483_G), .S(I_2482_S));
  generic_pmos I_2483(.D(I_2483_D), .G(I_2483_G), .S(I_2483_S));
  generic_nmos I_2484(.D(VSS), .G(I_2453_D), .S(I_2485_S));
  generic_pmos I_2485(.D(VDD), .G(I_2453_D), .S(I_2485_S));
  generic_nmos I_2486(.D(VSS), .G(I_2454_D), .S(I_2487_S));
  generic_pmos I_2487(.D(VDD), .G(I_2454_D), .S(I_2487_S));
  generic_nmos I_2488(.D(I_2489_D), .G(I_2425_D), .S(VSS));
  generic_pmos I_2489(.D(I_2489_D), .G(I_2425_D), .S(VDD));
  generic_pmos I_249(.D(I_281_D), .G(I_153_D), .S(VDD));
  generic_nmos I_2490(.D(I_2490_D), .G(I_2489_D), .S(I_2491_D));
  generic_pmos I_2491(.D(I_2491_D), .G(I_2489_D), .S(VDD));
  generic_nmos I_2492(.D(I_2492_D), .G(I_2650_D), .S(I_2493_D));
  generic_pmos I_2493(.D(I_2493_D), .G(I_2650_D), .S(VDD));
  generic_nmos I_2494(.D(I_2494_D), .G(I_2558_S), .S(VSS));
  generic_pmos I_2495(.D(I_2495_D), .G(I_2558_S), .S(VDD));
  generic_nmos I_2496(.D(I_2497_D), .G(I_2657_D), .S(I_2529_D));
  generic_pmos I_2497(.D(I_2497_D), .G(I_2625_S), .S(I_2529_D));
  generic_nmos I_2498(.D(I_2498_D), .G(I_2498_G), .S(VSS));
  generic_pmos I_2499(.D(I_2530_S), .G(I_2535_G), .S(VDD));
  generic_pmos I_25(.D(I_25_D), .G(I_25_G), .S(I_57_D));
  generic_nmos I_250(.D(VSS), .G(I_347_D), .S(I_251_S));
  generic_nmos I_2500(.D(I_2501_D), .G(I_2530_S), .S(I_2533_D));
  generic_pmos I_2501(.D(I_2501_D), .G(I_2535_G), .S(I_2533_D));
  generic_nmos I_2502(.D(I_2533_S), .G(I_2535_G), .S(I_2535_D));
  generic_pmos I_2503(.D(I_2533_S), .G(I_2534_G), .S(I_2535_D));
  generic_nmos I_2504(.D(I_2504_D), .G(I_2504_G), .S(I_2536_D));
  generic_pmos I_2505(.D(I_2505_D), .G(I_2536_G), .S(I_2537_D));
  generic_nmos I_2506(.D(VSS), .G(I_3751_S), .S(I_2539_S));
  generic_pmos I_2507(.D(VDD), .G(I_3591_S), .S(I_2539_D));
  generic_nmos I_2508(.D(VSS), .G(I_3591_S), .S(VSS));
  generic_pmos I_2509(.D(I_2509_D), .G(I_2540_G), .S(VDD));
  generic_pmos I_251(.D(VDD), .G(I_347_D), .S(I_251_S));
  generic_nmos I_2510(.D(I_2510_D), .G(I_2510_G), .S(I_2542_D));
  generic_pmos I_2511(.D(I_2511_D), .G(I_2542_G), .S(I_2543_D));
  generic_nmos I_2512(.D(I_3185_S), .G(I_2673_D), .S(I_2545_S));
  generic_pmos I_2513(.D(I_2513_D), .G(I_2544_G), .S(I_3185_S));
  generic_nmos I_2514(.D(I_2514_D), .G(I_2514_G), .S(I_2546_D));
  generic_pmos I_2515(.D(I_2515_D), .G(I_2546_G), .S(I_2547_D));
  generic_nmos I_2516(.D(I_2517_D), .G(I_2453_D), .S(I_2549_D));
  generic_pmos I_2517(.D(I_2517_D), .G(I_2485_S), .S(I_2549_D));
  generic_nmos I_2518(.D(VSS), .G(I_2454_D), .S(I_2869_D));
  generic_pmos I_2519(.D(I_2519_D), .G(I_2550_G), .S(I_2869_D));
  generic_nmos I_252(.D(VSS), .G(I_285_D), .S(I_253_S));
  generic_nmos I_2520(.D(I_2521_D), .G(I_1973_D), .S(I_2553_D));
  generic_pmos I_2521(.D(I_2521_D), .G(I_2007_D), .S(I_2553_D));
  generic_nmos I_2522(.D(VSS), .G(I_2427_D), .S(I_2554_D));
  generic_pmos I_2523(.D(VDD), .G(I_2871_D), .S(I_2555_D));
  generic_nmos I_2524(.D(VSS), .G(I_2429_D), .S(I_2556_D));
  generic_pmos I_2525(.D(VDD), .G(I_2653_D), .S(I_2557_D));
  generic_nmos I_2526(.D(I_2559_S), .G(I_2558_S), .S(VSS));
  generic_pmos I_2527(.D(I_2558_S), .G(I_1597_D), .S(VDD));
  generic_nmos I_2528(.D(I_2529_D), .G(I_2625_S), .S(I_2529_S));
  generic_pmos I_2529(.D(I_2529_D), .G(I_2657_D), .S(I_2529_S));
  generic_pmos I_253(.D(VDD), .G(I_285_D), .S(I_253_S));
  generic_nmos I_2530(.D(VSS), .G(I_2535_G), .S(I_2530_S));
  generic_pmos I_2531(.D(VDD), .G(I_2531_G), .S(I_2531_S));
  generic_nmos I_2532(.D(I_2533_D), .G(I_2535_G), .S(I_2533_S));
  generic_pmos I_2533(.D(I_2533_D), .G(I_2534_G), .S(I_2533_S));
  generic_nmos I_2534(.D(I_2535_D), .G(I_2534_G), .S(I_2535_S));
  generic_pmos I_2535(.D(I_2535_D), .G(I_2535_G), .S(I_2535_S));
  generic_nmos I_2536(.D(I_2536_D), .G(I_2536_G), .S(I_2536_S));
  generic_pmos I_2537(.D(I_2537_D), .G(I_2537_G), .S(I_2537_S));
  generic_nmos I_2538(.D(I_2539_S), .G(I_3591_S), .S(VSS));
  generic_pmos I_2539(.D(I_2539_D), .G(I_3751_S), .S(I_2539_S));
  generic_nmos I_254(.D(I_254_D), .G(I_255_G), .S(I_254_S));
  generic_nmos I_2540(.D(VSS), .G(I_2540_G), .S(I_2540_S));
  generic_pmos I_2541(.D(VDD), .G(I_3591_S), .S(VDD));
  generic_nmos I_2542(.D(I_2542_D), .G(I_2542_G), .S(I_2542_S));
  generic_pmos I_2543(.D(I_2543_D), .G(I_2543_G), .S(I_2543_S));
  generic_nmos I_2544(.D(I_2545_S), .G(I_2544_G), .S(I_2544_S));
  generic_pmos I_2545(.D(I_3185_S), .G(I_2705_S), .S(I_2545_S));
  generic_nmos I_2546(.D(I_2546_D), .G(I_2546_G), .S(I_2546_S));
  generic_pmos I_2547(.D(I_2547_D), .G(I_2547_G), .S(I_2547_S));
  generic_nmos I_2548(.D(I_2549_D), .G(I_2485_S), .S(I_2549_S));
  generic_pmos I_2549(.D(I_2549_D), .G(I_2453_D), .S(I_2549_S));
  generic_pmos I_255(.D(I_255_D), .G(I_255_G), .S(I_255_S));
  generic_nmos I_2550(.D(I_2869_D), .G(I_2550_G), .S(I_2550_S));
  generic_pmos I_2551(.D(I_2869_D), .G(I_2391_D), .S(VDD));
  generic_nmos I_2552(.D(I_2553_D), .G(I_2007_D), .S(I_2649_D));
  generic_pmos I_2553(.D(I_2553_D), .G(I_1973_D), .S(I_2649_D));
  generic_nmos I_2554(.D(I_2554_D), .G(I_2871_D), .S(I_2555_D));
  generic_pmos I_2555(.D(I_2555_D), .G(I_2427_D), .S(VDD));
  generic_nmos I_2556(.D(I_2556_D), .G(I_2653_D), .S(I_2557_D));
  generic_pmos I_2557(.D(I_2557_D), .G(I_2429_D), .S(VDD));
  generic_nmos I_2558(.D(VSS), .G(I_1597_D), .S(I_2558_S));
  generic_pmos I_2559(.D(VDD), .G(I_2558_S), .S(I_2559_S));
  generic_nmos I_256(.D(VSS), .G(I_227_D), .S(I_288_D));
  generic_nmos I_2560(.D(I_2657_D), .G(I_2561_G), .S(I_2592_D));
  generic_pmos I_2561(.D(VDD), .G(I_2561_G), .S(I_2657_D));
  generic_nmos I_2562(.D(I_2562_D), .G(I_2563_G), .S(I_2594_D));
  generic_pmos I_2563(.D(I_2563_D), .G(I_2563_G), .S(I_2595_D));
  generic_nmos I_2564(.D(I_2661_D), .G(I_2695_S), .S(VSS));
  generic_pmos I_2565(.D(I_2661_D), .G(I_2695_S), .S(VDD));
  generic_nmos I_2566(.D(I_2693_S), .G(I_2631_S), .S(I_2598_D));
  generic_pmos I_2567(.D(VDD), .G(I_2631_S), .S(I_2693_S));
  generic_nmos I_2568(.D(I_2632_D), .G(I_3493_S), .S(VSS));
  generic_pmos I_2569(.D(I_2632_D), .G(I_3493_S), .S(I_2601_D));
  generic_pmos I_257(.D(VDD), .G(I_1832_D), .S(I_289_D));
  generic_nmos I_2570(.D(I_2634_D), .G(I_3751_S), .S(VSS));
  generic_pmos I_2571(.D(I_2634_D), .G(I_3751_S), .S(I_2603_D));
  generic_nmos I_2572(.D(I_2572_D), .G(I_2573_G), .S(I_2604_D));
  generic_pmos I_2573(.D(I_2573_D), .G(I_2573_G), .S(I_2605_D));
  generic_nmos I_2574(.D(I_2574_D), .G(I_2575_G), .S(I_2606_D));
  generic_pmos I_2575(.D(I_2575_D), .G(I_2575_G), .S(I_2607_D));
  generic_nmos I_2576(.D(I_2576_D), .G(I_2577_G), .S(I_2609_D));
  generic_pmos I_2577(.D(I_2577_D), .G(I_2577_G), .S(I_2609_D));
  generic_nmos I_2578(.D(I_2578_D), .G(I_2579_G), .S(I_2610_D));
  generic_pmos I_2579(.D(I_2579_D), .G(I_2579_G), .S(I_2611_D));
  generic_nmos I_258(.D(I_291_D), .G(I_387_S), .S(I_290_D));
  generic_nmos I_2580(.D(I_2580_D), .G(I_2581_G), .S(I_2612_D));
  generic_pmos I_2581(.D(I_2581_D), .G(I_2581_G), .S(I_2613_D));
  generic_nmos I_2582(.D(I_2871_S), .G(I_2487_S), .S(I_2614_D));
  generic_pmos I_2583(.D(VDD), .G(I_2487_S), .S(I_2871_S));
  generic_nmos I_2584(.D(I_2585_D), .G(I_2553_D), .S(VSS));
  generic_pmos I_2585(.D(I_2585_D), .G(I_2553_D), .S(VDD));
  generic_nmos I_2586(.D(VSS), .G(I_2491_D), .S(I_2618_D));
  generic_pmos I_2587(.D(VDD), .G(I_2491_D), .S(I_2650_D));
  generic_nmos I_2588(.D(I_2653_D), .G(I_2495_D), .S(I_2620_D));
  generic_pmos I_2589(.D(I_2653_D), .G(I_2495_D), .S(VDD));
  generic_pmos I_259(.D(VDD), .G(I_549_S), .S(I_291_D));
  generic_nmos I_2590(.D(I_2655_D), .G(I_3593_S), .S(I_2622_D));
  generic_pmos I_2591(.D(I_2655_D), .G(I_3593_S), .S(VDD));
  generic_nmos I_2592(.D(I_2592_D), .G(I_2625_S), .S(VSS));
  generic_pmos I_2593(.D(I_2657_D), .G(I_2625_S), .S(VDD));
  generic_nmos I_2594(.D(I_2594_D), .G(I_2595_G), .S(I_2626_D));
  generic_pmos I_2595(.D(I_2595_D), .G(I_2595_G), .S(I_2627_D));
  generic_nmos I_2596(.D(VSS), .G(I_3241_D), .S(I_2628_D));
  generic_pmos I_2597(.D(VDD), .G(I_3241_D), .S(I_2695_S));
  generic_nmos I_2598(.D(I_2598_D), .G(I_3241_D), .S(VSS));
  generic_pmos I_2599(.D(I_2693_S), .G(I_3241_D), .S(VDD));
  generic_nmos I_26(.D(VSS), .G(I_1115_D), .S(I_59_D));
  generic_nmos I_260(.D(I_261_D), .G(I_329_D), .S(I_293_D));
  generic_nmos I_2600(.D(VSS), .G(I_3333_S), .S(I_2632_D));
  generic_pmos I_2601(.D(I_2601_D), .G(I_3333_S), .S(I_2633_D));
  generic_nmos I_2602(.D(VSS), .G(I_3493_S), .S(I_2634_D));
  generic_pmos I_2603(.D(I_2603_D), .G(I_3493_S), .S(I_2635_D));
  generic_nmos I_2604(.D(I_2604_D), .G(I_2605_G), .S(I_2636_D));
  generic_pmos I_2605(.D(I_2605_D), .G(I_2605_G), .S(I_2637_D));
  generic_nmos I_2606(.D(I_2606_D), .G(I_2607_G), .S(I_2638_D));
  generic_pmos I_2607(.D(I_2607_D), .G(I_2607_G), .S(I_2639_D));
  generic_nmos I_2608(.D(I_2609_D), .G(I_2545_S), .S(VSS));
  generic_pmos I_2609(.D(I_2609_D), .G(I_2545_S), .S(VDD));
  generic_pmos I_261(.D(I_261_D), .G(I_395_D), .S(I_293_D));
  generic_nmos I_2610(.D(I_2610_D), .G(I_2611_G), .S(I_2642_D));
  generic_pmos I_2611(.D(I_2611_D), .G(I_2611_G), .S(I_2643_D));
  generic_nmos I_2612(.D(I_2612_D), .G(I_2613_G), .S(I_2644_D));
  generic_pmos I_2613(.D(I_2613_D), .G(I_2613_G), .S(I_2645_D));
  generic_nmos I_2614(.D(I_2614_D), .G(I_2391_D), .S(VSS));
  generic_pmos I_2615(.D(I_2871_S), .G(I_2391_D), .S(VDD));
  generic_nmos I_2616(.D(VSS), .G(I_2585_D), .S(I_2649_D));
  generic_pmos I_2617(.D(VDD), .G(I_2585_D), .S(I_2649_D));
  generic_nmos I_2618(.D(I_2618_D), .G(I_2555_D), .S(I_2650_D));
  generic_pmos I_2619(.D(I_2650_D), .G(I_2555_D), .S(VDD));
  generic_nmos I_262(.D(I_263_D), .G(I_395_D), .S(I_295_D));
  generic_nmos I_2620(.D(I_2620_D), .G(I_2655_D), .S(I_2652_D));
  generic_pmos I_2621(.D(VDD), .G(I_2655_D), .S(I_2653_D));
  generic_nmos I_2622(.D(I_2622_D), .G(I_2558_S), .S(I_2654_D));
  generic_pmos I_2623(.D(VDD), .G(I_2558_S), .S(I_2655_D));
  generic_nmos I_2624(.D(VSS), .G(I_2689_D), .S(I_2625_S));
  generic_pmos I_2625(.D(VDD), .G(I_2689_D), .S(I_2625_S));
  generic_nmos I_2626(.D(I_2626_D), .G(I_2627_G), .S(I_2626_S));
  generic_pmos I_2627(.D(I_2627_D), .G(I_2627_G), .S(I_2627_S));
  generic_nmos I_2628(.D(I_2628_D), .G(I_2693_D), .S(I_2695_S));
  generic_pmos I_2629(.D(I_2695_S), .G(I_2693_D), .S(VDD));
  generic_pmos I_263(.D(I_263_D), .G(I_329_D), .S(I_295_D));
  generic_nmos I_2630(.D(VSS), .G(I_2695_D), .S(I_2631_S));
  generic_pmos I_2631(.D(VDD), .G(I_2695_D), .S(I_2631_S));
  generic_nmos I_2632(.D(I_2632_D), .G(I_3653_S), .S(VSS));
  generic_pmos I_2633(.D(I_2633_D), .G(I_3653_S), .S(VDD));
  generic_nmos I_2634(.D(I_2634_D), .G(I_3653_S), .S(VSS));
  generic_pmos I_2635(.D(I_2635_D), .G(I_3653_S), .S(VDD));
  generic_nmos I_2636(.D(I_2636_D), .G(I_2637_G), .S(I_2636_S));
  generic_pmos I_2637(.D(I_2637_D), .G(I_2637_G), .S(I_2637_S));
  generic_nmos I_2638(.D(I_2638_D), .G(I_2639_G), .S(I_2638_S));
  generic_pmos I_2639(.D(I_2639_D), .G(I_2639_G), .S(I_2639_S));
  generic_nmos I_264(.D(I_297_S), .G(I_616_S), .S(VSS));
  generic_nmos I_2640(.D(VSS), .G(I_2609_D), .S(I_2641_S));
  generic_pmos I_2641(.D(VDD), .G(I_2609_D), .S(I_2641_S));
  generic_nmos I_2642(.D(I_2642_D), .G(I_2643_G), .S(I_2642_S));
  generic_pmos I_2643(.D(I_2643_D), .G(I_2643_G), .S(I_2643_S));
  generic_nmos I_2644(.D(I_2644_D), .G(I_2645_G), .S(I_2644_S));
  generic_pmos I_2645(.D(I_2645_D), .G(I_2645_G), .S(I_2645_S));
  generic_nmos I_2646(.D(VSS), .G(I_2871_S), .S(I_2839_D));
  generic_pmos I_2647(.D(VDD), .G(I_2871_S), .S(I_2839_D));
  generic_nmos I_2648(.D(I_2649_D), .G(I_2585_D), .S(VSS));
  generic_pmos I_2649(.D(I_2649_D), .G(I_2585_D), .S(VDD));
  generic_pmos I_265(.D(I_265_D), .G(I_296_G), .S(VDD));
  generic_nmos I_2650(.D(I_2650_D), .G(I_2651_G), .S(I_2650_S));
  generic_pmos I_2651(.D(VDD), .G(I_2651_G), .S(I_2651_S));
  generic_nmos I_2652(.D(I_2652_D), .G(I_2815_D), .S(VSS));
  generic_pmos I_2653(.D(I_2653_D), .G(I_2815_D), .S(VDD));
  generic_nmos I_2654(.D(I_2654_D), .G(I_2719_S), .S(VSS));
  generic_pmos I_2655(.D(I_2655_D), .G(I_2719_S), .S(VDD));
  generic_nmos I_2656(.D(I_2657_D), .G(I_2945_S), .S(I_2689_D));
  generic_pmos I_2657(.D(I_2657_D), .G(I_3169_S), .S(I_2689_D));
  generic_nmos I_2658(.D(I_2658_D), .G(I_2658_G), .S(I_2690_D));
  generic_pmos I_2659(.D(I_2659_D), .G(I_2690_G), .S(I_2691_D));
  generic_nmos I_266(.D(I_266_D), .G(I_266_G), .S(I_298_D));
  generic_nmos I_2660(.D(I_2661_D), .G(I_2533_S), .S(I_2693_D));
  generic_pmos I_2661(.D(I_2661_D), .G(I_2471_S), .S(I_2693_D));
  generic_nmos I_2662(.D(I_2693_S), .G(I_2471_S), .S(I_2695_D));
  generic_pmos I_2663(.D(I_2693_S), .G(I_2533_S), .S(I_2695_D));
  generic_nmos I_2664(.D(I_2664_D), .G(I_2664_G), .S(I_2696_D));
  generic_pmos I_2665(.D(I_2665_D), .G(I_2696_G), .S(I_2697_D));
  generic_nmos I_2666(.D(I_2699_D), .G(I_2634_D), .S(I_2698_D));
  generic_pmos I_2667(.D(VDD), .G(I_2794_D), .S(I_2699_D));
  generic_nmos I_2668(.D(I_2668_D), .G(I_2668_G), .S(I_2700_D));
  generic_pmos I_2669(.D(I_2669_D), .G(I_2700_G), .S(I_2701_D));
  generic_pmos I_267(.D(I_267_D), .G(I_298_G), .S(I_299_D));
  generic_nmos I_2670(.D(I_3019_S), .G(I_2799_S), .S(I_3669_S));
  generic_pmos I_2671(.D(I_3019_S), .G(I_3823_S), .S(I_3669_S));
  generic_nmos I_2672(.D(I_2673_D), .G(I_2609_D), .S(I_3031_S));
  generic_pmos I_2673(.D(I_2673_D), .G(I_2641_S), .S(I_3031_S));
  generic_nmos I_2674(.D(I_2674_D), .G(I_2674_G), .S(I_2706_D));
  generic_pmos I_2675(.D(I_2675_D), .G(I_2706_G), .S(I_2707_D));
  generic_nmos I_2676(.D(I_2805_S), .G(I_2869_D), .S(I_2709_D));
  generic_pmos I_2677(.D(I_2805_S), .G(I_2741_D), .S(I_2709_D));
  generic_nmos I_2678(.D(I_2869_D), .G(I_2839_D), .S(I_2711_S));
  generic_pmos I_2679(.D(I_2679_D), .G(I_2710_G), .S(I_2869_D));
  generic_nmos I_268(.D(I_268_D), .G(I_268_G), .S(I_300_D));
  generic_nmos I_2680(.D(I_2681_D), .G(I_1973_D), .S(I_2713_D));
  generic_pmos I_2681(.D(I_2681_D), .G(I_2007_D), .S(I_2713_D));
  generic_nmos I_2682(.D(VSS), .G(I_2747_D), .S(I_2714_D));
  generic_pmos I_2683(.D(VDD), .G(I_2709_D), .S(I_2715_D));
  generic_nmos I_2684(.D(I_2717_D), .G(I_2493_D), .S(I_2716_D));
  generic_pmos I_2685(.D(VDD), .G(I_2557_D), .S(I_2717_D));
  generic_nmos I_2686(.D(I_2719_S), .G(I_2718_S), .S(VSS));
  generic_pmos I_2687(.D(I_2718_S), .G(I_1821_D), .S(VDD));
  generic_nmos I_2688(.D(I_2689_D), .G(I_3169_S), .S(I_2753_D));
  generic_pmos I_2689(.D(I_2689_D), .G(I_2945_S), .S(I_2753_D));
  generic_pmos I_269(.D(I_269_D), .G(I_300_G), .S(I_301_D));
  generic_nmos I_2690(.D(I_2690_D), .G(I_2690_G), .S(I_2690_S));
  generic_pmos I_2691(.D(I_2691_D), .G(I_2691_G), .S(I_2691_S));
  generic_nmos I_2692(.D(I_2693_D), .G(I_2471_S), .S(I_2693_S));
  generic_pmos I_2693(.D(I_2693_D), .G(I_2533_S), .S(I_2693_S));
  generic_nmos I_2694(.D(I_2695_D), .G(I_2533_S), .S(I_2695_S));
  generic_pmos I_2695(.D(I_2695_D), .G(I_2471_S), .S(I_2695_S));
  generic_nmos I_2696(.D(I_2696_D), .G(I_2696_G), .S(I_2696_S));
  generic_pmos I_2697(.D(I_2697_D), .G(I_2697_G), .S(I_2697_S));
  generic_nmos I_2698(.D(I_2698_D), .G(I_2794_D), .S(VSS));
  generic_pmos I_2699(.D(I_2699_D), .G(I_2634_D), .S(VDD));
  generic_pmos I_27(.D(VDD), .G(I_1115_D), .S(I_59_D));
  generic_nmos I_270(.D(I_270_D), .G(I_270_G), .S(I_302_D));
  generic_nmos I_2700(.D(I_2700_D), .G(I_2700_G), .S(I_2700_S));
  generic_pmos I_2701(.D(I_2701_D), .G(I_2701_G), .S(I_2701_S));
  generic_nmos I_2702(.D(I_3669_S), .G(I_3823_S), .S(I_2735_D));
  generic_pmos I_2703(.D(I_3669_S), .G(I_2799_S), .S(I_2735_D));
  generic_nmos I_2704(.D(I_3031_S), .G(I_2641_S), .S(I_2705_S));
  generic_pmos I_2705(.D(I_3031_S), .G(I_2609_D), .S(I_2705_S));
  generic_nmos I_2706(.D(I_2706_D), .G(I_2706_G), .S(I_2706_S));
  generic_pmos I_2707(.D(I_2707_D), .G(I_2707_G), .S(I_2707_S));
  generic_nmos I_2708(.D(I_2709_D), .G(I_2741_D), .S(I_2709_S));
  generic_pmos I_2709(.D(I_2709_D), .G(I_2869_D), .S(I_2709_S));
  generic_pmos I_271(.D(I_271_D), .G(I_302_G), .S(I_303_D));
  generic_nmos I_2710(.D(I_2711_S), .G(I_2710_G), .S(I_2710_S));
  generic_pmos I_2711(.D(I_2869_D), .G(I_2871_S), .S(I_2711_S));
  generic_nmos I_2712(.D(I_2713_D), .G(I_2007_D), .S(I_2809_D));
  generic_pmos I_2713(.D(I_2713_D), .G(I_1973_D), .S(I_2809_D));
  generic_nmos I_2714(.D(I_2714_D), .G(I_2709_D), .S(I_2715_D));
  generic_pmos I_2715(.D(I_2715_D), .G(I_2747_D), .S(VDD));
  generic_nmos I_2716(.D(I_2716_D), .G(I_2557_D), .S(VSS));
  generic_pmos I_2717(.D(I_2717_D), .G(I_2493_D), .S(VDD));
  generic_nmos I_2718(.D(VSS), .G(I_1821_D), .S(I_2718_S));
  generic_pmos I_2719(.D(VDD), .G(I_2718_S), .S(I_2719_S));
  generic_nmos I_272(.D(I_272_D), .G(I_272_G), .S(I_304_D));
  generic_nmos I_2720(.D(I_2753_D), .G(I_2849_D), .S(I_2752_D));
  generic_pmos I_2721(.D(VDD), .G(I_2849_D), .S(I_2753_D));
  generic_nmos I_2722(.D(I_2722_D), .G(I_2723_G), .S(I_2754_D));
  generic_pmos I_2723(.D(I_2723_D), .G(I_2723_G), .S(I_2755_D));
  generic_nmos I_2724(.D(I_2821_D), .G(I_2855_S), .S(VSS));
  generic_pmos I_2725(.D(I_2821_D), .G(I_2855_S), .S(VDD));
  generic_nmos I_2726(.D(I_2853_S), .G(I_2791_S), .S(I_2758_D));
  generic_pmos I_2727(.D(VDD), .G(I_2791_S), .S(I_2853_S));
  generic_nmos I_2728(.D(I_2728_D), .G(I_2729_G), .S(I_2760_D));
  generic_pmos I_2729(.D(I_2729_D), .G(I_2729_G), .S(I_2761_D));
  generic_pmos I_273(.D(I_273_D), .G(I_304_G), .S(I_305_D));
  generic_nmos I_2730(.D(I_2794_D), .G(I_2951_S), .S(VSS));
  generic_pmos I_2731(.D(I_2794_D), .G(I_2951_S), .S(I_2763_D));
  generic_nmos I_2732(.D(I_2732_D), .G(I_2733_G), .S(I_2764_D));
  generic_pmos I_2733(.D(I_2733_D), .G(I_2733_G), .S(I_2765_D));
  generic_nmos I_2734(.D(I_2735_D), .G(I_3019_S), .S(VSS));
  generic_pmos I_2735(.D(I_2735_D), .G(I_3019_S), .S(VDD));
  generic_nmos I_2736(.D(I_2736_D), .G(I_2737_G), .S(VSS));
  generic_pmos I_2737(.D(I_2737_D), .G(I_2737_G), .S(VDD));
  generic_nmos I_2738(.D(I_2738_D), .G(I_2739_G), .S(I_2770_D));
  generic_pmos I_2739(.D(I_2739_D), .G(I_2739_G), .S(I_2771_D));
  generic_nmos I_274(.D(I_274_D), .G(I_274_G), .S(I_306_D));
  generic_nmos I_2740(.D(I_2741_D), .G(I_2869_D), .S(VSS));
  generic_pmos I_2741(.D(I_2741_D), .G(I_2869_D), .S(VDD));
  generic_nmos I_2742(.D(I_2742_D), .G(I_2743_G), .S(I_2775_D));
  generic_pmos I_2743(.D(I_2743_D), .G(I_2743_G), .S(I_2775_D));
  generic_nmos I_2744(.D(I_2745_D), .G(I_2713_D), .S(VSS));
  generic_pmos I_2745(.D(I_2745_D), .G(I_2713_D), .S(VDD));
  generic_nmos I_2746(.D(I_2747_D), .G(I_1755_D), .S(VSS));
  generic_pmos I_2747(.D(I_2747_D), .G(I_1755_D), .S(VDD));
  generic_nmos I_2748(.D(I_2749_D), .G(I_2009_D), .S(VSS));
  generic_pmos I_2749(.D(I_2749_D), .G(I_2009_D), .S(VDD));
  generic_pmos I_275(.D(I_275_D), .G(I_306_G), .S(I_307_D));
  generic_nmos I_2750(.D(I_2815_D), .G(I_2559_S), .S(I_2782_D));
  generic_pmos I_2751(.D(I_2815_D), .G(I_2559_S), .S(VDD));
  generic_nmos I_2752(.D(I_2752_D), .G(I_2753_G), .S(VSS));
  generic_pmos I_2753(.D(I_2753_D), .G(I_2753_G), .S(VDD));
  generic_nmos I_2754(.D(I_2754_D), .G(I_2755_G), .S(I_2786_D));
  generic_pmos I_2755(.D(I_2755_D), .G(I_2755_G), .S(I_2787_D));
  generic_nmos I_2756(.D(VSS), .G(I_3241_D), .S(I_2788_D));
  generic_pmos I_2757(.D(VDD), .G(I_3241_D), .S(I_2855_S));
  generic_nmos I_2758(.D(I_2758_D), .G(I_3241_D), .S(VSS));
  generic_pmos I_2759(.D(I_2853_S), .G(I_3241_D), .S(VDD));
  generic_nmos I_276(.D(I_277_D), .G(I_341_D), .S(I_308_D));
  generic_nmos I_2760(.D(I_2760_D), .G(I_2761_G), .S(I_2792_D));
  generic_pmos I_2761(.D(I_2761_D), .G(I_2761_G), .S(I_2793_D));
  generic_nmos I_2762(.D(VSS), .G(I_3111_S), .S(I_2794_D));
  generic_pmos I_2763(.D(I_2763_D), .G(I_3111_S), .S(I_2795_D));
  generic_nmos I_2764(.D(I_2764_D), .G(I_2765_G), .S(I_2796_D));
  generic_pmos I_2765(.D(I_2765_D), .G(I_2765_G), .S(I_2797_D));
  generic_nmos I_2766(.D(VSS), .G(I_2767_G), .S(VSS));
  generic_pmos I_2767(.D(VDD), .G(I_2767_G), .S(VDD));
  generic_nmos I_2768(.D(VSS), .G(I_3065_D), .S(VSS));
  generic_pmos I_2769(.D(VDD), .G(I_3065_D), .S(VDD));
  generic_pmos I_277(.D(I_277_D), .G(I_341_D), .S(I_309_D));
  generic_nmos I_2770(.D(I_2770_D), .G(I_2771_G), .S(VSS));
  generic_pmos I_2771(.D(I_2771_D), .G(I_2771_G), .S(VDD));
  generic_nmos I_2772(.D(VSS), .G(I_2773_G), .S(VSS));
  generic_pmos I_2773(.D(VDD), .G(I_2773_G), .S(VDD));
  generic_nmos I_2774(.D(I_2775_D), .G(I_2711_S), .S(VSS));
  generic_pmos I_2775(.D(I_2775_D), .G(I_2711_S), .S(VDD));
  generic_nmos I_2776(.D(VSS), .G(I_2745_D), .S(I_2809_D));
  generic_pmos I_2777(.D(VDD), .G(I_2745_D), .S(I_2809_D));
  generic_nmos I_2778(.D(VSS), .G(I_1755_D), .S(I_2810_D));
  generic_pmos I_2779(.D(VDD), .G(I_1755_D), .S(I_2811_D));
  generic_nmos I_278(.D(I_279_D), .G(I_315_D), .S(I_311_D));
  generic_nmos I_2780(.D(VSS), .G(I_2009_D), .S(I_2812_D));
  generic_pmos I_2781(.D(VDD), .G(I_2009_D), .S(I_2813_D));
  generic_nmos I_2782(.D(I_2782_D), .G(I_2718_S), .S(I_2814_D));
  generic_pmos I_2783(.D(VDD), .G(I_2718_S), .S(I_2815_D));
  generic_nmos I_2784(.D(VSS), .G(I_2753_D), .S(I_2817_D));
  generic_pmos I_2785(.D(VDD), .G(I_2753_D), .S(I_2817_D));
  generic_nmos I_2786(.D(I_2786_D), .G(I_2787_G), .S(I_2786_S));
  generic_pmos I_2787(.D(I_2787_D), .G(I_2787_G), .S(I_2787_S));
  generic_nmos I_2788(.D(I_2788_D), .G(I_2853_D), .S(I_2855_S));
  generic_pmos I_2789(.D(I_2855_S), .G(I_2853_D), .S(VDD));
  generic_pmos I_279(.D(I_279_D), .G(I_251_S), .S(I_311_D));
  generic_nmos I_2790(.D(VSS), .G(I_2855_D), .S(I_2791_S));
  generic_pmos I_2791(.D(VDD), .G(I_2855_D), .S(I_2791_S));
  generic_nmos I_2792(.D(I_2792_D), .G(I_2793_G), .S(I_2792_S));
  generic_pmos I_2793(.D(I_2793_D), .G(I_2793_G), .S(I_2793_S));
  generic_nmos I_2794(.D(I_2794_D), .G(I_3271_S), .S(VSS));
  generic_pmos I_2795(.D(I_2795_D), .G(I_3271_S), .S(VDD));
  generic_nmos I_2796(.D(I_2796_D), .G(I_2797_G), .S(I_2796_S));
  generic_pmos I_2797(.D(I_2797_D), .G(I_2797_G), .S(I_2797_S));
  generic_nmos I_2798(.D(VSS), .G(I_3823_S), .S(I_2799_S));
  generic_pmos I_2799(.D(VDD), .G(I_3823_S), .S(I_2799_S));
  generic_nmos I_28(.D(VSS), .G(I_503_G), .S(I_93_S));
  generic_nmos I_280(.D(I_281_D), .G(I_251_S), .S(I_313_D));
  generic_nmos I_2800(.D(VSS), .G(I_2801_G), .S(I_2800_S));
  generic_pmos I_2801(.D(VDD), .G(I_2801_G), .S(I_2801_S));
  generic_nmos I_2802(.D(VSS), .G(I_2709_S), .S(VSS));
  generic_pmos I_2803(.D(VDD), .G(I_2709_S), .S(VDD));
  generic_nmos I_2804(.D(VSS), .G(I_2709_S), .S(I_2805_S));
  generic_pmos I_2805(.D(VDD), .G(I_2709_S), .S(I_2805_S));
  generic_nmos I_2806(.D(VSS), .G(I_2775_D), .S(I_2807_S));
  generic_pmos I_2807(.D(VDD), .G(I_2775_D), .S(I_2807_S));
  generic_nmos I_2808(.D(I_2809_D), .G(I_2745_D), .S(VSS));
  generic_pmos I_2809(.D(I_2809_D), .G(I_2745_D), .S(VDD));
  generic_pmos I_281(.D(I_281_D), .G(I_315_D), .S(I_313_D));
  generic_nmos I_2810(.D(I_2810_D), .G(I_2649_D), .S(I_2811_D));
  generic_pmos I_2811(.D(I_2811_D), .G(I_2649_D), .S(VDD));
  generic_nmos I_2812(.D(I_2812_D), .G(I_2875_D), .S(I_2813_D));
  generic_pmos I_2813(.D(I_2813_D), .G(I_2875_D), .S(VDD));
  generic_nmos I_2814(.D(I_2814_D), .G(I_2157_S), .S(VSS));
  generic_pmos I_2815(.D(I_2815_D), .G(I_2157_S), .S(VDD));
  generic_nmos I_2816(.D(I_2817_D), .G(I_3169_S), .S(I_2849_D));
  generic_pmos I_2817(.D(I_2817_D), .G(I_2945_S), .S(I_2849_D));
  generic_nmos I_2818(.D(I_2818_D), .G(I_2818_G), .S(I_2850_D));
  generic_pmos I_2819(.D(I_2819_D), .G(I_2850_G), .S(I_2851_D));
  generic_nmos I_282(.D(VSS), .G(I_251_S), .S(I_315_D));
  generic_nmos I_2820(.D(I_2821_D), .G(I_2693_S), .S(I_2853_D));
  generic_pmos I_2821(.D(I_2821_D), .G(I_2631_S), .S(I_2853_D));
  generic_nmos I_2822(.D(I_2853_S), .G(I_2631_S), .S(I_2855_D));
  generic_pmos I_2823(.D(I_2853_S), .G(I_2693_S), .S(I_2855_D));
  generic_nmos I_2824(.D(I_2824_D), .G(I_2824_G), .S(I_2856_D));
  generic_pmos I_2825(.D(I_2825_D), .G(I_2856_G), .S(I_2857_D));
  generic_nmos I_2826(.D(I_2826_D), .G(I_2826_G), .S(VSS));
  generic_pmos I_2827(.D(I_2955_D), .G(I_3751_S), .S(VDD));
  generic_nmos I_2828(.D(I_2828_D), .G(I_2828_G), .S(I_2860_D));
  generic_pmos I_2829(.D(I_2829_D), .G(I_2860_G), .S(I_2861_D));
  generic_pmos I_283(.D(VDD), .G(I_251_S), .S(I_315_D));
  generic_nmos I_2830(.D(I_2830_D), .G(I_2830_G), .S(I_2862_D));
  generic_pmos I_2831(.D(I_2831_D), .G(I_2862_G), .S(I_2863_D));
  generic_nmos I_2832(.D(I_2865_D), .G(I_1679_D), .S(I_2864_D));
  generic_pmos I_2833(.D(VDD), .G(I_3116_D), .S(I_2865_D));
  generic_nmos I_2834(.D(I_2834_D), .G(I_2834_G), .S(I_2866_D));
  generic_pmos I_2835(.D(I_2835_D), .G(I_2866_G), .S(I_2867_D));
  generic_nmos I_2836(.D(I_2869_D), .G(I_2709_S), .S(I_3191_D));
  generic_pmos I_2837(.D(I_2837_D), .G(I_2805_S), .S(I_2869_D));
  generic_nmos I_2838(.D(I_2839_D), .G(I_2775_D), .S(I_2871_D));
  generic_pmos I_2839(.D(I_2839_D), .G(I_2807_S), .S(I_2871_D));
  generic_nmos I_284(.D(I_285_D), .G(I_95_D), .S(I_317_D));
  generic_nmos I_2840(.D(I_2841_D), .G(I_1973_D), .S(I_2873_D));
  generic_pmos I_2841(.D(I_2841_D), .G(I_2007_D), .S(I_2873_D));
  generic_nmos I_2842(.D(I_2875_D), .G(I_2811_D), .S(I_2874_D));
  generic_pmos I_2843(.D(VDD), .G(I_2715_D), .S(I_2875_D));
  generic_nmos I_2844(.D(VSS), .G(I_2749_D), .S(I_2876_D));
  generic_pmos I_2845(.D(VDD), .G(I_3133_D), .S(I_2877_D));
  generic_nmos I_2846(.D(VSS), .G(I_2717_D), .S(I_2879_D));
  generic_pmos I_2847(.D(VDD), .G(I_2717_D), .S(I_2879_D));
  generic_nmos I_2848(.D(I_2849_D), .G(I_2945_S), .S(I_2849_S));
  generic_pmos I_2849(.D(I_2849_D), .G(I_3169_S), .S(I_2849_S));
  generic_pmos I_285(.D(I_285_D), .G(I_93_S), .S(I_317_D));
  generic_nmos I_2850(.D(I_2850_D), .G(I_2850_G), .S(I_2850_S));
  generic_pmos I_2851(.D(I_2851_D), .G(I_2851_G), .S(I_2851_S));
  generic_nmos I_2852(.D(I_2853_D), .G(I_2631_S), .S(I_2853_S));
  generic_pmos I_2853(.D(I_2853_D), .G(I_2693_S), .S(I_2853_S));
  generic_nmos I_2854(.D(I_2855_D), .G(I_2693_S), .S(I_2855_S));
  generic_pmos I_2855(.D(I_2855_D), .G(I_2631_S), .S(I_2855_S));
  generic_nmos I_2856(.D(I_2856_D), .G(I_2856_G), .S(I_2856_S));
  generic_pmos I_2857(.D(I_2857_D), .G(I_2857_G), .S(I_2857_S));
  generic_nmos I_2858(.D(VSS), .G(I_3751_S), .S(I_2890_D));
  generic_pmos I_2859(.D(VDD), .G(I_2859_G), .S(I_2859_S));
  generic_nmos I_286(.D(I_575_S), .G(I_93_S), .S(I_319_D));
  generic_nmos I_2860(.D(I_2860_D), .G(I_2860_G), .S(I_2860_S));
  generic_pmos I_2861(.D(I_2861_D), .G(I_2861_G), .S(I_2861_S));
  generic_nmos I_2862(.D(I_2862_D), .G(I_2862_G), .S(I_2862_S));
  generic_pmos I_2863(.D(I_2863_D), .G(I_2863_G), .S(I_2863_S));
  generic_nmos I_2864(.D(I_2864_D), .G(I_3116_D), .S(VSS));
  generic_pmos I_2865(.D(I_2865_D), .G(I_1679_D), .S(VDD));
  generic_nmos I_2866(.D(I_2866_D), .G(I_2866_G), .S(I_2866_S));
  generic_pmos I_2867(.D(I_2867_D), .G(I_2867_G), .S(I_2867_S));
  generic_nmos I_2868(.D(I_3191_D), .G(I_2805_S), .S(VSS));
  generic_pmos I_2869(.D(I_2869_D), .G(I_2805_S), .S(I_3191_D));
  generic_pmos I_287(.D(I_575_S), .G(I_95_D), .S(I_319_D));
  generic_nmos I_2870(.D(I_2871_D), .G(I_2807_S), .S(I_2871_S));
  generic_pmos I_2871(.D(I_2871_D), .G(I_2775_D), .S(I_2871_S));
  generic_nmos I_2872(.D(I_2873_D), .G(I_2007_D), .S(I_2969_D));
  generic_pmos I_2873(.D(I_2873_D), .G(I_1973_D), .S(I_2969_D));
  generic_nmos I_2874(.D(I_2874_D), .G(I_2715_D), .S(VSS));
  generic_pmos I_2875(.D(I_2875_D), .G(I_2811_D), .S(VDD));
  generic_nmos I_2876(.D(I_2876_D), .G(I_3133_D), .S(I_2877_D));
  generic_pmos I_2877(.D(I_2877_D), .G(I_2749_D), .S(VDD));
  generic_nmos I_2878(.D(I_2879_D), .G(I_2717_D), .S(VSS));
  generic_pmos I_2879(.D(I_2879_D), .G(I_2717_D), .S(VDD));
  generic_nmos I_288(.D(I_288_D), .G(I_1832_D), .S(I_289_D));
  generic_nmos I_2880(.D(I_3169_S), .G(I_2881_G), .S(I_2912_D));
  generic_pmos I_2881(.D(VDD), .G(I_2881_G), .S(I_3169_S));
  generic_nmos I_2882(.D(I_2882_D), .G(I_2883_G), .S(I_2914_D));
  generic_pmos I_2883(.D(I_2883_D), .G(I_2883_G), .S(I_2915_D));
  generic_nmos I_2884(.D(I_2981_D), .G(I_3015_S), .S(VSS));
  generic_pmos I_2885(.D(I_2981_D), .G(I_3015_S), .S(VDD));
  generic_nmos I_2886(.D(I_3013_S), .G(I_2951_S), .S(I_2918_D));
  generic_pmos I_2887(.D(VDD), .G(I_2951_S), .S(I_3013_S));
  generic_nmos I_2888(.D(I_2889_D), .G(I_1033_D), .S(VSS));
  generic_pmos I_2889(.D(I_2889_D), .G(I_1033_D), .S(VDD));
  generic_pmos I_289(.D(I_289_D), .G(I_227_D), .S(VDD));
  generic_nmos I_2890(.D(I_2890_D), .G(I_3271_S), .S(I_2922_D));
  generic_pmos I_2891(.D(I_2955_D), .G(I_3271_S), .S(VDD));
  generic_nmos I_2892(.D(I_2893_D), .G(I_2253_D), .S(VSS));
  generic_pmos I_2893(.D(I_2893_D), .G(I_2253_D), .S(VDD));
  generic_nmos I_2894(.D(I_2894_D), .G(I_2895_G), .S(VSS));
  generic_pmos I_2895(.D(I_2895_D), .G(I_2895_G), .S(VDD));
  generic_nmos I_2896(.D(VSS), .G(I_1679_D), .S(I_2928_D));
  generic_pmos I_2897(.D(I_2928_D), .G(I_1679_D), .S(I_2929_D));
  generic_nmos I_2898(.D(I_2898_D), .G(I_2899_G), .S(I_2930_D));
  generic_pmos I_2899(.D(I_2899_D), .G(I_2899_G), .S(I_2931_D));
  generic_pmos I_29(.D(VDD), .G(I_503_G), .S(I_93_S));
  generic_nmos I_290(.D(I_290_D), .G(I_549_S), .S(VSS));
  generic_nmos I_2900(.D(I_2900_D), .G(I_2901_G), .S(I_2932_D));
  generic_pmos I_2901(.D(I_2901_D), .G(I_2901_G), .S(I_2933_D));
  generic_nmos I_2902(.D(I_2902_D), .G(I_2903_G), .S(I_2934_D));
  generic_pmos I_2903(.D(I_2903_D), .G(I_2903_G), .S(I_2935_D));
  generic_nmos I_2904(.D(I_2905_D), .G(I_2873_D), .S(VSS));
  generic_pmos I_2905(.D(I_2905_D), .G(I_2873_D), .S(VDD));
  generic_nmos I_2906(.D(I_2907_D), .G(I_1755_D), .S(VSS));
  generic_pmos I_2907(.D(I_2907_D), .G(I_1755_D), .S(VDD));
  generic_nmos I_2908(.D(VSS), .G(I_2813_D), .S(I_2940_D));
  generic_pmos I_2909(.D(VDD), .G(I_2813_D), .S(I_2972_D));
  generic_pmos I_291(.D(I_291_D), .G(I_387_S), .S(VDD));
  generic_nmos I_2910(.D(I_2975_D), .G(I_3036_G), .S(I_2942_D));
  generic_pmos I_2911(.D(I_2975_D), .G(I_3036_G), .S(VDD));
  generic_nmos I_2912(.D(I_2912_D), .G(I_2945_S), .S(VSS));
  generic_pmos I_2913(.D(I_3169_S), .G(I_2945_S), .S(VDD));
  generic_nmos I_2914(.D(I_2914_D), .G(I_2915_G), .S(I_2946_D));
  generic_pmos I_2915(.D(I_2915_D), .G(I_2915_G), .S(I_2947_D));
  generic_nmos I_2916(.D(VSS), .G(I_3241_D), .S(I_2948_D));
  generic_pmos I_2917(.D(VDD), .G(I_3241_D), .S(I_3015_S));
  generic_nmos I_2918(.D(I_2918_D), .G(I_3241_D), .S(VSS));
  generic_pmos I_2919(.D(I_3013_S), .G(I_3241_D), .S(VDD));
  generic_nmos I_292(.D(I_293_D), .G(I_395_D), .S(I_293_S));
  generic_nmos I_2920(.D(VSS), .G(I_1033_D), .S(I_2952_D));
  generic_pmos I_2921(.D(VDD), .G(I_1033_D), .S(I_2953_D));
  generic_nmos I_2922(.D(I_2922_D), .G(I_2951_S), .S(I_2954_D));
  generic_pmos I_2923(.D(VDD), .G(I_2951_S), .S(I_2955_D));
  generic_nmos I_2924(.D(VSS), .G(I_2253_D), .S(I_2956_D));
  generic_pmos I_2925(.D(VDD), .G(I_2253_D), .S(I_2957_D));
  generic_nmos I_2926(.D(VSS), .G(I_3065_D), .S(VSS));
  generic_pmos I_2927(.D(VDD), .G(I_3065_D), .S(VDD));
  generic_nmos I_2928(.D(I_2928_D), .G(I_3116_D), .S(VSS));
  generic_pmos I_2929(.D(I_2929_D), .G(I_3116_D), .S(VDD));
  generic_pmos I_293(.D(I_293_D), .G(I_329_D), .S(I_293_S));
  generic_nmos I_2930(.D(I_2930_D), .G(I_2931_G), .S(I_2962_D));
  generic_pmos I_2931(.D(I_2931_D), .G(I_2931_G), .S(I_2963_D));
  generic_nmos I_2932(.D(I_2932_D), .G(I_2933_G), .S(I_2964_D));
  generic_pmos I_2933(.D(I_2933_D), .G(I_2933_G), .S(I_2965_D));
  generic_nmos I_2934(.D(I_2934_D), .G(I_2935_G), .S(I_2966_D));
  generic_pmos I_2935(.D(I_2935_D), .G(I_2935_G), .S(I_2967_D));
  generic_nmos I_2936(.D(VSS), .G(I_2905_D), .S(I_2969_D));
  generic_pmos I_2937(.D(VDD), .G(I_2905_D), .S(I_2969_D));
  generic_nmos I_2938(.D(VSS), .G(I_1755_D), .S(I_2970_D));
  generic_pmos I_2939(.D(VDD), .G(I_1755_D), .S(I_2971_D));
  generic_nmos I_294(.D(I_295_D), .G(I_329_D), .S(I_2329_D));
  generic_nmos I_2940(.D(I_2940_D), .G(I_2877_D), .S(I_2972_D));
  generic_pmos I_2941(.D(I_2972_D), .G(I_2877_D), .S(VDD));
  generic_nmos I_2942(.D(I_2942_D), .G(I_3198_S), .S(I_2974_D));
  generic_pmos I_2943(.D(VDD), .G(I_3198_S), .S(I_2975_D));
  generic_nmos I_2944(.D(VSS), .G(I_3009_D), .S(I_2945_S));
  generic_pmos I_2945(.D(VDD), .G(I_3009_D), .S(I_2945_S));
  generic_nmos I_2946(.D(I_2946_D), .G(I_2947_G), .S(I_2946_S));
  generic_pmos I_2947(.D(I_2947_D), .G(I_2947_G), .S(I_2947_S));
  generic_nmos I_2948(.D(I_2948_D), .G(I_3013_D), .S(I_3015_S));
  generic_pmos I_2949(.D(I_3015_S), .G(I_3013_D), .S(VDD));
  generic_pmos I_295(.D(I_295_D), .G(I_395_D), .S(I_2329_D));
  generic_nmos I_2950(.D(VSS), .G(I_3015_D), .S(I_2951_S));
  generic_pmos I_2951(.D(VDD), .G(I_3015_D), .S(I_2951_S));
  generic_nmos I_2952(.D(I_2952_D), .G(I_2955_D), .S(I_2953_D));
  generic_pmos I_2953(.D(I_2953_D), .G(I_2955_D), .S(VDD));
  generic_nmos I_2954(.D(I_2954_D), .G(I_3111_S), .S(I_2955_D));
  generic_pmos I_2955(.D(I_2955_D), .G(I_3111_S), .S(VDD));
  generic_nmos I_2956(.D(I_2956_D), .G(I_3339_D), .S(I_2957_D));
  generic_pmos I_2957(.D(I_2957_D), .G(I_3339_D), .S(VDD));
  generic_nmos I_2958(.D(VSS), .G(I_2959_G), .S(I_2958_S));
  generic_pmos I_2959(.D(VDD), .G(I_2959_G), .S(I_2959_S));
  generic_nmos I_296(.D(VSS), .G(I_296_G), .S(I_296_S));
  generic_nmos I_2960(.D(VSS), .G(I_2928_D), .S(I_2961_S));
  generic_pmos I_2961(.D(VDD), .G(I_2928_D), .S(I_2961_S));
  generic_nmos I_2962(.D(I_2962_D), .G(I_2963_G), .S(I_2962_S));
  generic_pmos I_2963(.D(I_2963_D), .G(I_2963_G), .S(I_2963_S));
  generic_nmos I_2964(.D(I_2964_D), .G(I_2965_G), .S(I_2964_S));
  generic_pmos I_2965(.D(I_2965_D), .G(I_2965_G), .S(I_2965_S));
  generic_nmos I_2966(.D(I_2966_D), .G(I_2967_G), .S(I_2966_S));
  generic_pmos I_2967(.D(I_2967_D), .G(I_2967_G), .S(I_2967_S));
  generic_nmos I_2968(.D(I_2969_D), .G(I_2905_D), .S(VSS));
  generic_pmos I_2969(.D(I_2969_D), .G(I_2905_D), .S(VDD));
  generic_pmos I_297(.D(VDD), .G(I_616_S), .S(I_297_S));
  generic_nmos I_2970(.D(I_2970_D), .G(I_2809_D), .S(I_2971_D));
  generic_pmos I_2971(.D(I_2971_D), .G(I_2809_D), .S(VDD));
  generic_nmos I_2972(.D(I_2972_D), .G(I_2973_G), .S(I_2972_S));
  generic_pmos I_2973(.D(VDD), .G(I_2973_G), .S(I_2973_S));
  generic_nmos I_2974(.D(I_2974_D), .G(I_3038_S), .S(VSS));
  generic_pmos I_2975(.D(I_2975_D), .G(I_3038_S), .S(VDD));
  generic_nmos I_2976(.D(I_3169_S), .G(I_3265_S), .S(I_3009_D));
  generic_pmos I_2977(.D(I_3169_S), .G(I_3489_S), .S(I_3009_D));
  generic_nmos I_2978(.D(I_3075_D), .G(I_2632_D), .S(I_3010_D));
  generic_pmos I_2979(.D(VDD), .G(I_2791_S), .S(I_3075_D));
  generic_nmos I_298(.D(I_298_D), .G(I_298_G), .S(I_298_S));
  generic_nmos I_2980(.D(I_2981_D), .G(I_2853_S), .S(I_3013_D));
  generic_pmos I_2981(.D(I_2981_D), .G(I_2791_S), .S(I_3013_D));
  generic_nmos I_2982(.D(I_3013_S), .G(I_2791_S), .S(I_3015_D));
  generic_pmos I_2983(.D(I_3013_S), .G(I_2853_S), .S(I_3015_D));
  generic_nmos I_2984(.D(VSS), .G(I_2889_D), .S(I_3016_D));
  generic_pmos I_2985(.D(VDD), .G(I_3083_D), .S(I_3017_D));
  generic_nmos I_2986(.D(I_3019_S), .G(I_3019_G), .S(VSS));
  generic_pmos I_2987(.D(I_2987_D), .G(I_3018_G), .S(VDD));
  generic_nmos I_2988(.D(VSS), .G(I_2893_D), .S(I_3020_D));
  generic_pmos I_2989(.D(VDD), .G(I_3271_S), .S(I_3021_D));
  generic_pmos I_299(.D(I_299_D), .G(I_299_G), .S(I_299_S));
  generic_nmos I_2990(.D(I_3023_D), .G(I_3116_D), .S(I_3022_D));
  generic_pmos I_2991(.D(VDD), .G(I_3019_S), .S(I_3023_D));
  generic_nmos I_2992(.D(VSS), .G(I_2928_D), .S(I_3825_S));
  generic_pmos I_2993(.D(I_2993_D), .G(I_3024_G), .S(I_3825_S));
  generic_nmos I_2994(.D(I_3123_S), .G(I_3219_D), .S(I_3027_D));
  generic_pmos I_2995(.D(I_3123_S), .G(I_3059_D), .S(I_3027_D));
  generic_nmos I_2996(.D(I_3125_S), .G(I_3191_S), .S(I_3029_D));
  generic_pmos I_2997(.D(I_3125_S), .G(I_3061_D), .S(I_3029_D));
  generic_nmos I_2998(.D(I_3127_S), .G(I_3191_D), .S(I_3031_D));
  generic_pmos I_2999(.D(I_3127_S), .G(I_3063_D), .S(I_3031_D));
  generic_pmos I_3(.D(I_3_D), .G(I_3_G), .S(VDD));
  generic_nmos I_30(.D(I_95_D), .G(I_95_G), .S(VSS));
  generic_nmos I_300(.D(I_300_D), .G(I_300_G), .S(I_300_S));
  generic_nmos I_3000(.D(I_3993_S), .G(I_1973_D), .S(I_3033_D));
  generic_pmos I_3001(.D(I_3993_S), .G(I_2007_D), .S(I_3033_D));
  generic_nmos I_3002(.D(VSS), .G(I_2907_D), .S(I_3034_D));
  generic_pmos I_3003(.D(VDD), .G(I_3031_D), .S(I_3035_D));
  generic_nmos I_3004(.D(I_3004_D), .G(I_3004_G), .S(VSS));
  generic_pmos I_3005(.D(I_3036_S), .G(I_3036_G), .S(VDD));
  generic_nmos I_3006(.D(I_3039_S), .G(I_3038_S), .S(VSS));
  generic_pmos I_3007(.D(I_3038_S), .G(I_1597_D), .S(VDD));
  generic_nmos I_3008(.D(I_3009_D), .G(I_3489_S), .S(I_3073_D));
  generic_pmos I_3009(.D(I_3009_D), .G(I_3265_S), .S(I_3073_D));
  generic_pmos I_301(.D(I_301_D), .G(I_301_G), .S(I_301_S));
  generic_nmos I_3010(.D(I_3010_D), .G(I_2791_S), .S(I_3042_D));
  generic_pmos I_3011(.D(I_3075_D), .G(I_2632_D), .S(VDD));
  generic_nmos I_3012(.D(I_3013_D), .G(I_2791_S), .S(I_3013_S));
  generic_pmos I_3013(.D(I_3013_D), .G(I_2853_S), .S(I_3013_S));
  generic_nmos I_3014(.D(I_3015_D), .G(I_2853_S), .S(I_3015_S));
  generic_pmos I_3015(.D(I_3015_D), .G(I_2791_S), .S(I_3015_S));
  generic_nmos I_3016(.D(I_3016_D), .G(I_3083_D), .S(I_3017_D));
  generic_pmos I_3017(.D(I_3017_D), .G(I_2889_D), .S(VDD));
  generic_nmos I_3018(.D(VSS), .G(I_3018_G), .S(I_3018_S));
  generic_pmos I_3019(.D(VDD), .G(I_3019_G), .S(I_3019_S));
  generic_nmos I_302(.D(I_302_D), .G(I_302_G), .S(I_302_S));
  generic_nmos I_3020(.D(I_3020_D), .G(I_3271_S), .S(I_3021_D));
  generic_pmos I_3021(.D(I_3021_D), .G(I_2893_D), .S(VDD));
  generic_nmos I_3022(.D(I_3022_D), .G(I_3019_S), .S(VSS));
  generic_pmos I_3023(.D(I_3023_D), .G(I_3116_D), .S(VDD));
  generic_nmos I_3024(.D(I_3825_S), .G(I_3024_G), .S(I_3024_S));
  generic_pmos I_3025(.D(I_3825_S), .G(I_2865_D), .S(VDD));
  generic_nmos I_3026(.D(I_3027_D), .G(I_3059_D), .S(I_3985_D));
  generic_pmos I_3027(.D(I_3027_D), .G(I_3219_D), .S(I_3985_D));
  generic_nmos I_3028(.D(I_3029_D), .G(I_3061_D), .S(I_3345_D));
  generic_pmos I_3029(.D(I_3029_D), .G(I_3191_S), .S(I_3345_D));
  generic_pmos I_303(.D(I_303_D), .G(I_303_G), .S(I_303_S));
  generic_nmos I_3030(.D(I_3031_D), .G(I_3063_D), .S(I_3031_S));
  generic_pmos I_3031(.D(I_3031_D), .G(I_3191_D), .S(I_3031_S));
  generic_nmos I_3032(.D(I_3033_D), .G(I_2007_D), .S(I_3129_D));
  generic_pmos I_3033(.D(I_3033_D), .G(I_1973_D), .S(I_3129_D));
  generic_nmos I_3034(.D(I_3034_D), .G(I_3031_D), .S(I_3035_D));
  generic_pmos I_3035(.D(I_3035_D), .G(I_2907_D), .S(VDD));
  generic_nmos I_3036(.D(VSS), .G(I_3036_G), .S(I_3036_S));
  generic_pmos I_3037(.D(VDD), .G(I_3037_G), .S(I_3037_S));
  generic_nmos I_3038(.D(VSS), .G(I_1597_D), .S(I_3038_S));
  generic_pmos I_3039(.D(VDD), .G(I_3038_S), .S(I_3039_S));
  generic_nmos I_304(.D(I_304_D), .G(I_304_G), .S(I_304_S));
  generic_nmos I_3040(.D(I_3073_D), .G(I_3169_D), .S(I_3072_D));
  generic_pmos I_3041(.D(VDD), .G(I_3169_D), .S(I_3073_D));
  generic_nmos I_3042(.D(I_3042_D), .G(I_3173_S), .S(I_3074_D));
  generic_pmos I_3043(.D(VDD), .G(I_3173_S), .S(I_3075_D));
  generic_nmos I_3044(.D(I_3141_D), .G(I_3175_S), .S(VSS));
  generic_pmos I_3045(.D(I_3141_D), .G(I_3175_S), .S(VDD));
  generic_nmos I_3046(.D(I_3173_S), .G(I_3111_S), .S(I_3078_D));
  generic_pmos I_3047(.D(VDD), .G(I_3111_S), .S(I_3173_S));
  generic_nmos I_3048(.D(VSS), .G(I_2953_D), .S(I_3080_D));
  generic_pmos I_3049(.D(VDD), .G(I_2953_D), .S(I_3112_D));
  generic_pmos I_305(.D(I_305_D), .G(I_305_G), .S(I_305_S));
  generic_nmos I_3050(.D(I_3083_D), .G(I_2951_S), .S(I_3082_D));
  generic_pmos I_3051(.D(VDD), .G(I_2951_S), .S(I_3083_D));
  generic_nmos I_3052(.D(VSS), .G(I_2957_D), .S(I_3084_D));
  generic_pmos I_3053(.D(VDD), .G(I_2957_D), .S(I_3116_D));
  generic_nmos I_3054(.D(VSS), .G(I_3116_D), .S(I_3086_D));
  generic_pmos I_3055(.D(I_3086_D), .G(I_3116_D), .S(I_3087_D));
  generic_nmos I_3056(.D(I_3345_S), .G(I_2961_S), .S(I_3088_D));
  generic_pmos I_3057(.D(VDD), .G(I_2961_S), .S(I_3345_S));
  generic_nmos I_3058(.D(I_3059_D), .G(I_3219_D), .S(VSS));
  generic_pmos I_3059(.D(I_3059_D), .G(I_3219_D), .S(VDD));
  generic_nmos I_306(.D(I_306_D), .G(I_306_G), .S(I_306_S));
  generic_nmos I_3060(.D(I_3061_D), .G(I_3191_S), .S(VSS));
  generic_pmos I_3061(.D(I_3061_D), .G(I_3191_S), .S(VDD));
  generic_nmos I_3062(.D(I_3063_D), .G(I_3191_D), .S(VSS));
  generic_pmos I_3063(.D(I_3063_D), .G(I_3191_D), .S(VDD));
  generic_nmos I_3064(.D(I_3065_D), .G(I_3033_D), .S(VSS));
  generic_pmos I_3065(.D(I_3065_D), .G(I_3033_D), .S(VDD));
  generic_nmos I_3066(.D(VSS), .G(I_2971_D), .S(I_3098_D));
  generic_pmos I_3067(.D(VDD), .G(I_2971_D), .S(I_3130_D));
  generic_nmos I_3068(.D(I_3133_D), .G(I_2975_D), .S(I_3100_D));
  generic_pmos I_3069(.D(I_3133_D), .G(I_2975_D), .S(VDD));
  generic_pmos I_307(.D(I_307_D), .G(I_307_G), .S(I_307_S));
  generic_nmos I_3070(.D(I_3135_D), .G(I_3659_S), .S(I_3102_D));
  generic_pmos I_3071(.D(I_3135_D), .G(I_3659_S), .S(VDD));
  generic_nmos I_3072(.D(I_3072_D), .G(I_3073_G), .S(VSS));
  generic_pmos I_3073(.D(I_3073_D), .G(I_3073_G), .S(VDD));
  generic_nmos I_3074(.D(I_3074_D), .G(I_3171_D), .S(VSS));
  generic_pmos I_3075(.D(I_3075_D), .G(I_3171_D), .S(VDD));
  generic_nmos I_3076(.D(VSS), .G(I_3241_D), .S(I_3108_D));
  generic_pmos I_3077(.D(VDD), .G(I_3241_D), .S(I_3175_S));
  generic_nmos I_3078(.D(I_3078_D), .G(I_3241_D), .S(VSS));
  generic_pmos I_3079(.D(I_3173_S), .G(I_3241_D), .S(VDD));
  generic_nmos I_308(.D(I_308_D), .G(I_341_D), .S(VSS));
  generic_nmos I_3080(.D(I_3080_D), .G(I_3017_D), .S(I_3112_D));
  generic_pmos I_3081(.D(I_3112_D), .G(I_3017_D), .S(VDD));
  generic_nmos I_3082(.D(I_3082_D), .G(I_3657_D), .S(VSS));
  generic_pmos I_3083(.D(I_3083_D), .G(I_3657_D), .S(VDD));
  generic_nmos I_3084(.D(I_3084_D), .G(I_3021_D), .S(I_3116_D));
  generic_pmos I_3085(.D(I_3116_D), .G(I_3021_D), .S(VDD));
  generic_nmos I_3086(.D(I_3086_D), .G(I_3019_S), .S(VSS));
  generic_pmos I_3087(.D(I_3087_D), .G(I_3019_S), .S(VDD));
  generic_nmos I_3088(.D(I_3088_D), .G(I_2865_D), .S(VSS));
  generic_pmos I_3089(.D(I_3345_S), .G(I_2865_D), .S(VDD));
  generic_pmos I_309(.D(I_309_D), .G(I_341_D), .S(VDD));
  generic_nmos I_3090(.D(VSS), .G(I_3091_G), .S(VSS));
  generic_pmos I_3091(.D(VDD), .G(I_3091_G), .S(VDD));
  generic_nmos I_3092(.D(VSS), .G(I_3093_G), .S(VSS));
  generic_pmos I_3093(.D(VDD), .G(I_3093_G), .S(VDD));
  generic_nmos I_3094(.D(VSS), .G(I_3095_G), .S(VSS));
  generic_pmos I_3095(.D(VDD), .G(I_3095_G), .S(VDD));
  generic_nmos I_3096(.D(VSS), .G(I_3065_D), .S(I_3129_D));
  generic_pmos I_3097(.D(VDD), .G(I_3065_D), .S(I_3129_D));
  generic_nmos I_3098(.D(I_3098_D), .G(I_3035_D), .S(I_3130_D));
  generic_pmos I_3099(.D(I_3130_D), .G(I_3035_D), .S(VDD));
  generic_pmos I_31(.D(I_95_D), .G(I_95_G), .S(VDD));
  generic_nmos I_310(.D(I_311_D), .G(I_251_S), .S(I_375_D));
  generic_nmos I_3100(.D(I_3100_D), .G(I_3135_D), .S(I_3132_D));
  generic_pmos I_3101(.D(VDD), .G(I_3135_D), .S(I_3133_D));
  generic_nmos I_3102(.D(I_3102_D), .G(I_3038_S), .S(I_3134_D));
  generic_pmos I_3103(.D(VDD), .G(I_3038_S), .S(I_3135_D));
  generic_nmos I_3104(.D(VSS), .G(I_3073_D), .S(I_3137_D));
  generic_pmos I_3105(.D(VDD), .G(I_3073_D), .S(I_3137_D));
  generic_nmos I_3106(.D(VSS), .G(I_3107_G), .S(I_3106_S));
  generic_pmos I_3107(.D(VDD), .G(I_3107_G), .S(I_3107_S));
  generic_nmos I_3108(.D(I_3108_D), .G(I_3173_D), .S(I_3175_S));
  generic_pmos I_3109(.D(I_3175_S), .G(I_3173_D), .S(VDD));
  generic_pmos I_311(.D(I_311_D), .G(I_315_D), .S(I_375_D));
  generic_nmos I_3110(.D(VSS), .G(I_3175_D), .S(I_3111_S));
  generic_pmos I_3111(.D(VDD), .G(I_3175_D), .S(I_3111_S));
  generic_nmos I_3112(.D(I_3112_D), .G(I_3113_G), .S(I_3112_S));
  generic_pmos I_3113(.D(VDD), .G(I_3113_G), .S(I_3113_S));
  generic_nmos I_3114(.D(VSS), .G(I_3115_G), .S(I_3114_S));
  generic_pmos I_3115(.D(VDD), .G(I_3115_G), .S(I_3115_S));
  generic_nmos I_3116(.D(I_3116_D), .G(I_3117_G), .S(I_3116_S));
  generic_pmos I_3117(.D(VDD), .G(I_3117_G), .S(I_3117_S));
  generic_nmos I_3118(.D(VSS), .G(I_3086_D), .S(I_3119_S));
  generic_pmos I_3119(.D(VDD), .G(I_3086_D), .S(I_3119_S));
  generic_nmos I_312(.D(I_313_D), .G(I_315_D), .S(I_409_S));
  generic_nmos I_3120(.D(VSS), .G(I_3345_S), .S(I_3313_D));
  generic_pmos I_3121(.D(VDD), .G(I_3345_S), .S(I_3313_D));
  generic_nmos I_3122(.D(VSS), .G(I_3985_D), .S(I_3123_S));
  generic_pmos I_3123(.D(VDD), .G(I_3985_D), .S(I_3123_S));
  generic_nmos I_3124(.D(VSS), .G(I_3345_D), .S(I_3125_S));
  generic_pmos I_3125(.D(VDD), .G(I_3345_D), .S(I_3125_S));
  generic_nmos I_3126(.D(VSS), .G(I_3031_S), .S(I_3127_S));
  generic_pmos I_3127(.D(VDD), .G(I_3031_S), .S(I_3127_S));
  generic_nmos I_3128(.D(I_3129_D), .G(I_3065_D), .S(VSS));
  generic_pmos I_3129(.D(I_3129_D), .G(I_3065_D), .S(VDD));
  generic_pmos I_313(.D(I_313_D), .G(I_251_S), .S(I_409_S));
  generic_nmos I_3130(.D(I_3130_D), .G(I_3131_G), .S(I_3130_S));
  generic_pmos I_3131(.D(VDD), .G(I_3131_G), .S(I_3131_S));
  generic_nmos I_3132(.D(I_3132_D), .G(I_3295_D), .S(VSS));
  generic_pmos I_3133(.D(I_3133_D), .G(I_3295_D), .S(VDD));
  generic_nmos I_3134(.D(I_3134_D), .G(I_3199_S), .S(VSS));
  generic_pmos I_3135(.D(I_3135_D), .G(I_3199_S), .S(VDD));
  generic_nmos I_3136(.D(I_3137_D), .G(I_3489_S), .S(I_3169_D));
  generic_pmos I_3137(.D(I_3137_D), .G(I_3265_S), .S(I_3169_D));
  generic_nmos I_3138(.D(I_3171_D), .G(I_3173_S), .S(I_3170_D));
  generic_pmos I_3139(.D(VDD), .G(I_3013_S), .S(I_3171_D));
  generic_nmos I_314(.D(I_315_D), .G(I_251_S), .S(VSS));
  generic_nmos I_3140(.D(I_3141_D), .G(I_3013_S), .S(I_3173_D));
  generic_pmos I_3141(.D(I_3141_D), .G(I_2951_S), .S(I_3173_D));
  generic_nmos I_3142(.D(I_3173_S), .G(I_2951_S), .S(I_3175_D));
  generic_pmos I_3143(.D(I_3173_S), .G(I_3013_S), .S(I_3175_D));
  generic_nmos I_3144(.D(VSS), .G(I_3112_D), .S(I_3176_D));
  generic_pmos I_3145(.D(VDD), .G(I_1283_D), .S(I_3177_D));
  generic_nmos I_3146(.D(I_3146_D), .G(I_3146_G), .S(I_3178_D));
  generic_pmos I_3147(.D(I_3147_D), .G(I_3178_G), .S(I_3179_D));
  generic_nmos I_3148(.D(I_3148_D), .G(I_3148_G), .S(I_3180_D));
  generic_pmos I_3149(.D(I_3149_D), .G(I_3593_S), .S(I_3181_D));
  generic_pmos I_315(.D(I_315_D), .G(I_251_S), .S(VDD));
  generic_nmos I_3150(.D(VSS), .G(I_3086_D), .S(I_3823_D));
  generic_pmos I_3151(.D(I_3151_D), .G(I_3182_G), .S(I_3823_D));
  generic_nmos I_3152(.D(I_3825_S), .G(I_3313_D), .S(I_3185_S));
  generic_pmos I_3153(.D(I_3153_D), .G(I_3184_G), .S(I_3825_S));
  generic_nmos I_3154(.D(I_3219_D), .G(I_3985_D), .S(I_3507_D));
  generic_pmos I_3155(.D(I_3155_D), .G(I_3123_S), .S(I_3219_D));
  generic_nmos I_3156(.D(I_3191_S), .G(I_3345_D), .S(I_3189_S));
  generic_pmos I_3157(.D(I_3157_D), .G(I_3125_S), .S(I_3191_S));
  generic_nmos I_3158(.D(I_3191_D), .G(I_3031_S), .S(I_3191_S));
  generic_pmos I_3159(.D(I_3159_D), .G(I_3127_S), .S(I_3191_D));
  generic_nmos I_316(.D(I_317_D), .G(I_93_S), .S(I_445_D));
  generic_nmos I_3160(.D(VSS), .G(I_3225_D), .S(I_3192_D));
  generic_pmos I_3161(.D(VDD), .G(I_3449_D), .S(I_3193_D));
  generic_nmos I_3162(.D(I_3195_S), .G(I_3195_G), .S(VSS));
  generic_pmos I_3163(.D(I_3163_D), .G(I_3194_G), .S(VDD));
  generic_nmos I_3164(.D(VSS), .G(I_3229_D), .S(I_3196_D));
  generic_pmos I_3165(.D(VDD), .G(I_3453_D), .S(I_3197_D));
  generic_nmos I_3166(.D(I_3199_S), .G(I_3198_S), .S(VSS));
  generic_pmos I_3167(.D(I_3198_S), .G(I_1821_D), .S(VDD));
  generic_nmos I_3168(.D(I_3169_D), .G(I_3265_S), .S(I_3169_S));
  generic_pmos I_3169(.D(I_3169_D), .G(I_3489_S), .S(I_3169_S));
  generic_pmos I_317(.D(I_317_D), .G(I_95_D), .S(I_445_D));
  generic_nmos I_3170(.D(I_3170_D), .G(I_3013_S), .S(VSS));
  generic_pmos I_3171(.D(I_3171_D), .G(I_3173_S), .S(VDD));
  generic_nmos I_3172(.D(I_3173_D), .G(I_2951_S), .S(I_3173_S));
  generic_pmos I_3173(.D(I_3173_D), .G(I_3013_S), .S(I_3173_S));
  generic_nmos I_3174(.D(I_3175_D), .G(I_3013_S), .S(I_3175_S));
  generic_pmos I_3175(.D(I_3175_D), .G(I_2951_S), .S(I_3175_S));
  generic_nmos I_3176(.D(I_3176_D), .G(I_1283_D), .S(I_3177_D));
  generic_pmos I_3177(.D(I_3177_D), .G(I_3112_D), .S(VDD));
  generic_nmos I_3178(.D(I_3178_D), .G(I_3178_G), .S(I_3178_S));
  generic_pmos I_3179(.D(I_3179_D), .G(I_3179_G), .S(I_3179_S));
  generic_nmos I_318(.D(I_319_D), .G(I_95_D), .S(I_415_S));
  generic_nmos I_3180(.D(I_3180_D), .G(I_3593_S), .S(I_3180_S));
  generic_pmos I_3181(.D(I_3181_D), .G(I_3181_G), .S(I_3181_S));
  generic_nmos I_3182(.D(I_3823_D), .G(I_3182_G), .S(I_3182_S));
  generic_pmos I_3183(.D(I_3823_D), .G(I_3023_D), .S(VDD));
  generic_nmos I_3184(.D(I_3185_S), .G(I_3184_G), .S(I_3184_S));
  generic_pmos I_3185(.D(I_3825_S), .G(I_3345_S), .S(I_3185_S));
  generic_nmos I_3186(.D(I_3507_D), .G(I_3123_S), .S(VSS));
  generic_pmos I_3187(.D(I_3219_D), .G(I_3123_S), .S(I_3507_D));
  generic_nmos I_3188(.D(I_3189_S), .G(I_3125_S), .S(VSS));
  generic_pmos I_3189(.D(I_3191_S), .G(I_3125_S), .S(I_3189_S));
  generic_pmos I_319(.D(I_319_D), .G(I_93_S), .S(I_415_S));
  generic_nmos I_3190(.D(I_3191_S), .G(I_3127_S), .S(VSS));
  generic_pmos I_3191(.D(I_3191_D), .G(I_3127_S), .S(I_3191_S));
  generic_nmos I_3192(.D(I_3192_D), .G(I_3449_D), .S(I_3193_D));
  generic_pmos I_3193(.D(I_3193_D), .G(I_3225_D), .S(VDD));
  generic_nmos I_3194(.D(VSS), .G(I_3194_G), .S(I_3194_S));
  generic_pmos I_3195(.D(VDD), .G(I_3195_G), .S(I_3195_S));
  generic_nmos I_3196(.D(I_3196_D), .G(I_3453_D), .S(I_3197_D));
  generic_pmos I_3197(.D(I_3197_D), .G(I_3229_D), .S(VDD));
  generic_nmos I_3198(.D(VSS), .G(I_1821_D), .S(I_3198_S));
  generic_pmos I_3199(.D(VDD), .G(I_3198_S), .S(I_3199_S));
  generic_nmos I_32(.D(I_32_D), .G(I_65_S), .S(VSS));
  generic_nmos I_320(.D(I_321_D), .G(I_33_D), .S(VSS));
  generic_nmos I_3200(.D(I_3489_S), .G(I_3201_G), .S(I_3232_D));
  generic_pmos I_3201(.D(VDD), .G(I_3201_G), .S(I_3489_S));
  generic_nmos I_3202(.D(I_3202_D), .G(I_3203_G), .S(I_3234_D));
  generic_pmos I_3203(.D(I_3203_D), .G(I_3203_G), .S(I_3235_D));
  generic_nmos I_3204(.D(I_3301_D), .G(I_3335_S), .S(VSS));
  generic_pmos I_3205(.D(I_3301_D), .G(I_3335_S), .S(VDD));
  generic_nmos I_3206(.D(I_3333_S), .G(I_3271_S), .S(I_3238_D));
  generic_pmos I_3207(.D(VDD), .G(I_3271_S), .S(I_3333_S));
  generic_nmos I_3208(.D(VSS), .G(I_3177_D), .S(I_3241_D));
  generic_pmos I_3209(.D(VDD), .G(I_3177_D), .S(I_3241_D));
  generic_pmos I_321(.D(I_321_D), .G(I_33_D), .S(VDD));
  generic_nmos I_3210(.D(I_3210_D), .G(I_3211_G), .S(I_3242_D));
  generic_pmos I_3211(.D(I_3211_D), .G(I_3211_G), .S(I_3243_D));
  generic_nmos I_3212(.D(I_3212_D), .G(I_3213_G), .S(I_3244_D));
  generic_pmos I_3213(.D(I_3213_D), .G(I_3213_G), .S(I_3245_D));
  generic_nmos I_3214(.D(I_3503_S), .G(I_3119_S), .S(I_3246_D));
  generic_pmos I_3215(.D(VDD), .G(I_3119_S), .S(I_3503_S));
  generic_nmos I_3216(.D(I_3216_D), .G(I_3217_G), .S(I_3249_D));
  generic_pmos I_3217(.D(I_3217_D), .G(I_3217_G), .S(I_3249_D));
  generic_nmos I_3218(.D(I_3219_D), .G(I_3283_S), .S(VSS));
  generic_pmos I_3219(.D(I_3219_D), .G(I_3283_S), .S(VDD));
  generic_nmos I_322(.D(I_355_D), .G(I_1029_D), .S(I_354_D));
  generic_nmos I_3220(.D(I_3220_D), .G(I_3221_G), .S(VSS));
  generic_pmos I_3221(.D(I_3221_D), .G(I_3221_G), .S(VDD));
  generic_nmos I_3222(.D(I_3287_D), .G(I_3347_D), .S(I_3254_D));
  generic_pmos I_3223(.D(I_3287_D), .G(I_3347_D), .S(VDD));
  generic_nmos I_3224(.D(I_3225_D), .G(I_1689_D), .S(VSS));
  generic_pmos I_3225(.D(I_3225_D), .G(I_1689_D), .S(VDD));
  generic_nmos I_3226(.D(I_3291_D), .G(VDD), .S(I_3258_D));
  generic_pmos I_3227(.D(I_3291_D), .G(VDD), .S(VDD));
  generic_nmos I_3228(.D(I_3229_D), .G(I_2009_D), .S(VSS));
  generic_pmos I_3229(.D(I_3229_D), .G(I_2009_D), .S(VDD));
  generic_pmos I_323(.D(VDD), .G(I_1029_D), .S(I_355_D));
  generic_nmos I_3230(.D(I_3295_D), .G(I_3039_S), .S(I_3262_D));
  generic_pmos I_3231(.D(I_3295_D), .G(I_3039_S), .S(VDD));
  generic_nmos I_3232(.D(I_3232_D), .G(I_3265_S), .S(VSS));
  generic_pmos I_3233(.D(I_3489_S), .G(I_3265_S), .S(VDD));
  generic_nmos I_3234(.D(I_3234_D), .G(I_3235_G), .S(I_3266_D));
  generic_pmos I_3235(.D(I_3235_D), .G(I_3235_G), .S(I_3267_D));
  generic_nmos I_3236(.D(VSS), .G(I_3241_D), .S(I_3268_D));
  generic_pmos I_3237(.D(VDD), .G(I_3241_D), .S(I_3335_S));
  generic_nmos I_3238(.D(I_3238_D), .G(I_3241_D), .S(VSS));
  generic_pmos I_3239(.D(I_3333_S), .G(I_3241_D), .S(VDD));
  generic_nmos I_324(.D(I_421_D), .G(I_1187_S), .S(I_356_D));
  generic_nmos I_3240(.D(I_3241_D), .G(I_3177_D), .S(VSS));
  generic_pmos I_3241(.D(I_3241_D), .G(I_3177_D), .S(VDD));
  generic_nmos I_3242(.D(I_3242_D), .G(I_3243_G), .S(VSS));
  generic_pmos I_3243(.D(I_3243_D), .G(I_3243_G), .S(VDD));
  generic_nmos I_3244(.D(I_3244_D), .G(I_3245_G), .S(I_3276_D));
  generic_pmos I_3245(.D(I_3245_D), .G(I_3245_G), .S(I_3277_D));
  generic_nmos I_3246(.D(I_3246_D), .G(I_3023_D), .S(VSS));
  generic_pmos I_3247(.D(I_3503_S), .G(I_3023_D), .S(VDD));
  generic_nmos I_3248(.D(I_3249_D), .G(I_3185_S), .S(VSS));
  generic_pmos I_3249(.D(I_3249_D), .G(I_3185_S), .S(VDD));
  generic_pmos I_325(.D(VDD), .G(I_1187_S), .S(I_421_D));
  generic_nmos I_3250(.D(VSS), .G(I_3251_G), .S(VSS));
  generic_pmos I_3251(.D(VDD), .G(I_3251_G), .S(VDD));
  generic_nmos I_3252(.D(VSS), .G(I_3349_D), .S(I_3284_D));
  generic_pmos I_3253(.D(VDD), .G(I_3349_D), .S(I_3285_D));
  generic_nmos I_3254(.D(I_3254_D), .G(I_3510_S), .S(I_3286_D));
  generic_pmos I_3255(.D(VDD), .G(I_3510_S), .S(I_3287_D));
  generic_nmos I_3256(.D(VSS), .G(I_1689_D), .S(I_3288_D));
  generic_pmos I_3257(.D(VDD), .G(I_1689_D), .S(I_3289_D));
  generic_nmos I_3258(.D(I_3258_D), .G(I_3514_S), .S(I_3290_D));
  generic_pmos I_3259(.D(VDD), .G(I_3514_S), .S(I_3291_D));
  generic_nmos I_326(.D(I_423_D), .G(I_453_S), .S(VSS));
  generic_nmos I_3260(.D(VSS), .G(I_2009_D), .S(I_3292_D));
  generic_pmos I_3261(.D(VDD), .G(I_2009_D), .S(I_3293_D));
  generic_nmos I_3262(.D(I_3262_D), .G(I_3198_S), .S(I_3294_D));
  generic_pmos I_3263(.D(VDD), .G(I_3198_S), .S(I_3295_D));
  generic_nmos I_3264(.D(VSS), .G(I_3329_D), .S(I_3265_S));
  generic_pmos I_3265(.D(VDD), .G(I_3329_D), .S(I_3265_S));
  generic_nmos I_3266(.D(I_3266_D), .G(I_3267_G), .S(I_3266_S));
  generic_pmos I_3267(.D(I_3267_D), .G(I_3267_G), .S(I_3267_S));
  generic_nmos I_3268(.D(I_3268_D), .G(I_3333_D), .S(I_3335_S));
  generic_pmos I_3269(.D(I_3335_S), .G(I_3333_D), .S(VDD));
  generic_pmos I_327(.D(I_423_D), .G(I_453_S), .S(VDD));
  generic_nmos I_3270(.D(VSS), .G(I_3335_D), .S(I_3271_S));
  generic_pmos I_3271(.D(VDD), .G(I_3335_D), .S(I_3271_S));
  generic_nmos I_3272(.D(VSS), .G(I_3591_S), .S(VSS));
  generic_pmos I_3273(.D(VDD), .G(I_3591_S), .S(VDD));
  generic_nmos I_3274(.D(VSS), .G(I_3591_S), .S(VSS));
  generic_pmos I_3275(.D(VDD), .G(I_3591_S), .S(VDD));
  generic_nmos I_3276(.D(I_3276_D), .G(I_3277_G), .S(I_3276_S));
  generic_pmos I_3277(.D(I_3277_D), .G(I_3277_G), .S(I_3277_S));
  generic_nmos I_3278(.D(VSS), .G(I_3503_S), .S(I_3471_D));
  generic_pmos I_3279(.D(VDD), .G(I_3503_S), .S(I_3471_D));
  generic_nmos I_328(.D(I_329_D), .G(I_395_D), .S(VSS));
  generic_nmos I_3280(.D(VSS), .G(I_3249_D), .S(I_3281_S));
  generic_pmos I_3281(.D(VDD), .G(I_3249_D), .S(I_3281_S));
  generic_nmos I_3282(.D(VSS), .G(I_3189_S), .S(I_3283_S));
  generic_pmos I_3283(.D(VDD), .G(I_3189_S), .S(I_3283_S));
  generic_nmos I_3284(.D(I_3284_D), .G(I_3413_D), .S(I_3285_D));
  generic_pmos I_3285(.D(I_3285_D), .G(I_3413_D), .S(VDD));
  generic_nmos I_3286(.D(I_3286_D), .G(I_3350_S), .S(VSS));
  generic_pmos I_3287(.D(I_3287_D), .G(I_3350_S), .S(VDD));
  generic_nmos I_3288(.D(I_3288_D), .G(I_3285_D), .S(I_3289_D));
  generic_pmos I_3289(.D(I_3289_D), .G(I_3285_D), .S(VDD));
  generic_pmos I_329(.D(I_329_D), .G(I_395_D), .S(VDD));
  generic_nmos I_3290(.D(I_3290_D), .G(I_3354_S), .S(VSS));
  generic_pmos I_3291(.D(I_3291_D), .G(I_3354_S), .S(VDD));
  generic_nmos I_3292(.D(I_3292_D), .G(I_3130_D), .S(I_3293_D));
  generic_pmos I_3293(.D(I_3293_D), .G(I_3130_D), .S(VDD));
  generic_nmos I_3294(.D(I_3294_D), .G(VSS), .S(VSS));
  generic_pmos I_3295(.D(I_3295_D), .G(VSS), .S(VDD));
  generic_nmos I_3296(.D(I_3489_S), .G(I_3555_G), .S(I_3329_D));
  generic_pmos I_3297(.D(I_3489_S), .G(I_3521_D), .S(I_3329_D));
  generic_nmos I_3298(.D(VSS), .G(I_3331_G), .S(I_3331_D));
  generic_pmos I_3299(.D(VDD), .G(I_3331_G), .S(I_3331_D));
  generic_pmos I_33(.D(I_33_D), .G(I_65_S), .S(VDD));
  generic_nmos I_330(.D(I_395_D), .G(I_618_S), .S(I_362_D));
  generic_nmos I_3300(.D(I_3301_D), .G(I_3173_S), .S(I_3333_D));
  generic_pmos I_3301(.D(I_3301_D), .G(I_3111_S), .S(I_3333_D));
  generic_nmos I_3302(.D(I_3333_S), .G(I_3111_S), .S(I_3335_D));
  generic_pmos I_3303(.D(I_3333_S), .G(I_3173_S), .S(I_3335_D));
  generic_nmos I_3304(.D(I_3433_S), .G(I_3591_S), .S(I_3337_D));
  generic_pmos I_3305(.D(I_3433_S), .G(I_3369_D), .S(I_3337_D));
  generic_nmos I_3306(.D(I_3435_S), .G(I_3499_D), .S(I_3339_D));
  generic_pmos I_3307(.D(I_3435_S), .G(I_3371_D), .S(I_3339_D));
  generic_nmos I_3308(.D(I_3308_D), .G(I_3308_G), .S(I_3340_D));
  generic_pmos I_3309(.D(I_3309_D), .G(I_3340_G), .S(I_3341_D));
  generic_pmos I_331(.D(I_395_D), .G(I_618_S), .S(VDD));
  generic_nmos I_3310(.D(I_3823_D), .G(I_3471_D), .S(I_3535_D));
  generic_pmos I_3311(.D(I_3311_D), .G(I_3342_G), .S(I_3823_D));
  generic_nmos I_3312(.D(I_3313_D), .G(I_3249_D), .S(I_3345_D));
  generic_pmos I_3313(.D(I_3313_D), .G(I_3281_S), .S(I_3345_D));
  generic_nmos I_3314(.D(I_3443_S), .G(I_3507_D), .S(I_3347_D));
  generic_pmos I_3315(.D(I_3443_S), .G(I_3379_D), .S(I_3347_D));
  generic_nmos I_3316(.D(I_3349_D), .G(I_3445_S), .S(I_3348_D));
  generic_pmos I_3317(.D(VDD), .G(I_1831_S), .S(I_3349_D));
  generic_nmos I_3318(.D(I_3351_S), .G(I_3350_S), .S(VSS));
  generic_pmos I_3319(.D(I_3350_S), .G(I_1597_D), .S(VDD));
  generic_nmos I_332(.D(I_332_D), .G(I_333_G), .S(I_364_D));
  generic_nmos I_3320(.D(I_3353_D), .G(I_3289_D), .S(I_3352_D));
  generic_pmos I_3321(.D(VDD), .G(I_3193_D), .S(I_3353_D));
  generic_nmos I_3322(.D(I_3355_S), .G(I_3354_S), .S(VSS));
  generic_pmos I_3323(.D(I_3354_S), .G(I_1597_D), .S(VDD));
  generic_nmos I_3324(.D(I_3357_D), .G(I_3293_D), .S(I_3356_D));
  generic_pmos I_3325(.D(VDD), .G(I_3197_D), .S(I_3357_D));
  generic_nmos I_3326(.D(VSS), .G(I_2972_D), .S(I_3359_D));
  generic_pmos I_3327(.D(VDD), .G(I_2972_D), .S(I_3359_D));
  generic_nmos I_3328(.D(I_3329_D), .G(I_3521_D), .S(I_3393_D));
  generic_pmos I_3329(.D(I_3329_D), .G(I_3555_G), .S(I_3393_D));
  generic_pmos I_333(.D(I_333_D), .G(I_333_G), .S(I_365_D));
  generic_nmos I_3330(.D(I_3331_D), .G(I_3331_G), .S(VSS));
  generic_pmos I_3331(.D(I_3331_D), .G(I_3331_G), .S(VDD));
  generic_nmos I_3332(.D(I_3333_D), .G(I_3111_S), .S(I_3333_S));
  generic_pmos I_3333(.D(I_3333_D), .G(I_3173_S), .S(I_3333_S));
  generic_nmos I_3334(.D(I_3335_D), .G(I_3173_S), .S(I_3335_S));
  generic_pmos I_3335(.D(I_3335_D), .G(I_3111_S), .S(I_3335_S));
  generic_nmos I_3336(.D(I_3337_D), .G(I_3369_D), .S(I_3499_D));
  generic_pmos I_3337(.D(I_3337_D), .G(I_3591_S), .S(I_3499_D));
  generic_nmos I_3338(.D(I_3339_D), .G(I_3371_D), .S(I_3497_S));
  generic_pmos I_3339(.D(I_3339_D), .G(I_3499_D), .S(I_3497_S));
  generic_nmos I_334(.D(I_334_D), .G(I_335_G), .S(I_366_D));
  generic_nmos I_3340(.D(I_3340_D), .G(I_3340_G), .S(I_3340_S));
  generic_pmos I_3341(.D(I_3341_D), .G(I_3341_G), .S(I_3341_S));
  generic_nmos I_3342(.D(I_3535_D), .G(I_3342_G), .S(I_3342_S));
  generic_pmos I_3343(.D(I_3823_D), .G(I_3503_S), .S(I_3535_D));
  generic_nmos I_3344(.D(I_3345_D), .G(I_3281_S), .S(I_3345_S));
  generic_pmos I_3345(.D(I_3345_D), .G(I_3249_D), .S(I_3345_S));
  generic_nmos I_3346(.D(I_3347_D), .G(I_3379_D), .S(I_3503_D));
  generic_pmos I_3347(.D(I_3347_D), .G(I_3507_D), .S(I_3503_D));
  generic_nmos I_3348(.D(I_3348_D), .G(I_1831_S), .S(VSS));
  generic_pmos I_3349(.D(I_3349_D), .G(I_3445_S), .S(VDD));
  generic_pmos I_335(.D(I_335_D), .G(I_335_G), .S(I_367_D));
  generic_nmos I_3350(.D(VSS), .G(I_1597_D), .S(I_3350_S));
  generic_pmos I_3351(.D(VDD), .G(I_3350_S), .S(I_3351_S));
  generic_nmos I_3352(.D(I_3352_D), .G(I_3193_D), .S(VSS));
  generic_pmos I_3353(.D(I_3353_D), .G(I_3289_D), .S(VDD));
  generic_nmos I_3354(.D(VSS), .G(I_1597_D), .S(I_3354_S));
  generic_pmos I_3355(.D(VDD), .G(I_3354_S), .S(I_3355_S));
  generic_nmos I_3356(.D(I_3356_D), .G(I_3197_D), .S(VSS));
  generic_pmos I_3357(.D(I_3357_D), .G(I_3293_D), .S(VDD));
  generic_nmos I_3358(.D(I_3359_D), .G(I_2972_D), .S(VSS));
  generic_pmos I_3359(.D(I_3359_D), .G(I_2972_D), .S(VDD));
  generic_nmos I_336(.D(I_336_D), .G(I_337_G), .S(I_368_D));
  generic_nmos I_3360(.D(I_3393_D), .G(I_3489_D), .S(I_3392_D));
  generic_pmos I_3361(.D(VDD), .G(I_3489_D), .S(I_3393_D));
  generic_nmos I_3362(.D(I_3363_D), .G(I_3491_S), .S(VSS));
  generic_pmos I_3363(.D(I_3363_D), .G(I_3491_S), .S(VDD));
  generic_nmos I_3364(.D(I_3461_D), .G(I_3495_S), .S(VSS));
  generic_pmos I_3365(.D(I_3461_D), .G(I_3495_S), .S(VDD));
  generic_nmos I_3366(.D(I_3493_S), .G(I_3431_S), .S(I_3398_D));
  generic_pmos I_3367(.D(VDD), .G(I_3431_S), .S(I_3493_S));
  generic_nmos I_3368(.D(I_3369_D), .G(I_3591_S), .S(VSS));
  generic_pmos I_3369(.D(I_3369_D), .G(I_3591_S), .S(VDD));
  generic_pmos I_337(.D(I_337_D), .G(I_337_G), .S(I_369_D));
  generic_nmos I_3370(.D(I_3371_D), .G(I_3499_D), .S(VSS));
  generic_pmos I_3371(.D(I_3371_D), .G(I_3499_D), .S(VDD));
  generic_nmos I_3372(.D(VSS), .G(I_3659_S), .S(VSS));
  generic_pmos I_3373(.D(VDD), .G(I_3659_S), .S(VDD));
  generic_nmos I_3374(.D(I_3374_D), .G(I_3375_G), .S(I_3407_D));
  generic_pmos I_3375(.D(I_3375_D), .G(I_3375_G), .S(I_3407_D));
  generic_nmos I_3376(.D(I_3376_D), .G(I_3377_G), .S(I_3408_D));
  generic_pmos I_3377(.D(I_3377_D), .G(I_3377_G), .S(I_3409_D));
  generic_nmos I_3378(.D(I_3379_D), .G(I_3507_D), .S(VSS));
  generic_pmos I_3379(.D(I_3379_D), .G(I_3507_D), .S(VDD));
  generic_nmos I_338(.D(I_338_D), .G(I_339_G), .S(I_370_D));
  generic_nmos I_3380(.D(I_3413_D), .G(I_3381_G), .S(I_3412_D));
  generic_pmos I_3381(.D(VDD), .G(I_3381_G), .S(I_3413_D));
  generic_nmos I_3382(.D(I_3447_D), .G(I_3987_S), .S(I_3414_D));
  generic_pmos I_3383(.D(I_3447_D), .G(I_3987_S), .S(VDD));
  generic_nmos I_3384(.D(I_3449_D), .G(I_3287_D), .S(I_3416_D));
  generic_pmos I_3385(.D(I_3449_D), .G(I_3287_D), .S(VDD));
  generic_nmos I_3386(.D(I_3451_D), .G(I_3983_D), .S(I_3418_D));
  generic_pmos I_3387(.D(I_3451_D), .G(I_3983_D), .S(VDD));
  generic_nmos I_3388(.D(I_3453_D), .G(I_3291_D), .S(I_3420_D));
  generic_pmos I_3389(.D(I_3453_D), .G(I_3291_D), .S(VDD));
  generic_pmos I_339(.D(I_339_D), .G(I_339_G), .S(I_371_D));
  generic_nmos I_3390(.D(VSS), .G(I_3357_D), .S(I_3423_D));
  generic_pmos I_3391(.D(VDD), .G(I_3357_D), .S(I_3423_D));
  generic_nmos I_3392(.D(I_3392_D), .G(I_3393_G), .S(VSS));
  generic_pmos I_3393(.D(I_3393_D), .G(I_3393_G), .S(VDD));
  generic_nmos I_3394(.D(VSS), .G(I_2853_S), .S(I_3426_D));
  generic_pmos I_3395(.D(VDD), .G(I_2853_S), .S(I_3427_D));
  generic_nmos I_3396(.D(VSS), .G(I_3241_D), .S(I_3428_D));
  generic_pmos I_3397(.D(VDD), .G(I_3241_D), .S(I_3495_S));
  generic_nmos I_3398(.D(I_3398_D), .G(I_3241_D), .S(VSS));
  generic_pmos I_3399(.D(I_3493_S), .G(I_3241_D), .S(VDD));
  generic_nmos I_34(.D(VSS), .G(I_3_D), .S(I_67_S));
  generic_nmos I_340(.D(I_341_D), .G(I_437_D), .S(I_372_D));
  generic_nmos I_3400(.D(VSS), .G(I_3401_G), .S(VSS));
  generic_pmos I_3401(.D(VDD), .G(I_3401_G), .S(VDD));
  generic_nmos I_3402(.D(VSS), .G(I_3403_G), .S(VSS));
  generic_pmos I_3403(.D(VDD), .G(I_3403_G), .S(VDD));
  generic_nmos I_3404(.D(VSS), .G(I_3501_D), .S(I_3436_D));
  generic_pmos I_3405(.D(VDD), .G(I_3501_D), .S(I_3663_S));
  generic_nmos I_3406(.D(I_3407_D), .G(I_3535_D), .S(VSS));
  generic_pmos I_3407(.D(I_3407_D), .G(I_3535_D), .S(VDD));
  generic_nmos I_3408(.D(I_3408_D), .G(I_3409_G), .S(I_3440_D));
  generic_pmos I_3409(.D(I_3409_D), .G(I_3409_G), .S(I_3441_D));
  generic_pmos I_341(.D(I_341_D), .G(I_437_D), .S(I_373_D));
  generic_nmos I_3410(.D(VSS), .G(I_3411_G), .S(VSS));
  generic_pmos I_3411(.D(VDD), .G(I_3411_G), .S(VDD));
  generic_nmos I_3412(.D(I_3412_D), .G(I_3735_G), .S(VSS));
  generic_pmos I_3413(.D(I_3413_D), .G(I_3735_G), .S(VDD));
  generic_nmos I_3414(.D(I_3414_D), .G(I_3350_S), .S(I_3446_D));
  generic_pmos I_3415(.D(VDD), .G(I_3350_S), .S(I_3447_D));
  generic_nmos I_3416(.D(I_3416_D), .G(I_3447_D), .S(I_3448_D));
  generic_pmos I_3417(.D(VDD), .G(I_3447_D), .S(I_3449_D));
  generic_nmos I_3418(.D(I_3418_D), .G(I_3354_S), .S(I_3450_D));
  generic_pmos I_3419(.D(VDD), .G(I_3354_S), .S(I_3451_D));
  generic_nmos I_342(.D(VSS), .G(I_471_D), .S(I_375_D));
  generic_nmos I_3420(.D(I_3420_D), .G(I_3451_D), .S(I_3452_D));
  generic_pmos I_3421(.D(VDD), .G(I_3451_D), .S(I_3453_D));
  generic_nmos I_3422(.D(I_3423_D), .G(I_3357_D), .S(VSS));
  generic_pmos I_3423(.D(I_3423_D), .G(I_3357_D), .S(VDD));
  generic_nmos I_3424(.D(VSS), .G(I_3393_D), .S(I_3457_D));
  generic_pmos I_3425(.D(VDD), .G(I_3393_D), .S(I_3457_D));
  generic_nmos I_3426(.D(I_3426_D), .G(I_3013_S), .S(I_3427_D));
  generic_pmos I_3427(.D(I_3427_D), .G(I_3013_S), .S(VDD));
  generic_nmos I_3428(.D(I_3428_D), .G(I_3493_D), .S(I_3495_S));
  generic_pmos I_3429(.D(I_3495_S), .G(I_3493_D), .S(VDD));
  generic_pmos I_343(.D(VDD), .G(I_471_D), .S(I_375_D));
  generic_nmos I_3430(.D(VSS), .G(I_3495_D), .S(I_3431_S));
  generic_pmos I_3431(.D(VDD), .G(I_3495_D), .S(I_3431_S));
  generic_nmos I_3432(.D(VSS), .G(I_3499_D), .S(I_3433_S));
  generic_pmos I_3433(.D(VDD), .G(I_3499_D), .S(I_3433_S));
  generic_nmos I_3434(.D(VSS), .G(I_3497_S), .S(I_3435_S));
  generic_pmos I_3435(.D(VDD), .G(I_3497_S), .S(I_3435_S));
  generic_nmos I_3436(.D(I_3436_D), .G(I_3565_D), .S(I_3663_S));
  generic_pmos I_3437(.D(I_3663_S), .G(I_3565_D), .S(VDD));
  generic_nmos I_3438(.D(VSS), .G(I_3407_D), .S(I_3439_S));
  generic_pmos I_3439(.D(VDD), .G(I_3407_D), .S(I_3439_S));
  generic_nmos I_344(.D(VSS), .G(I_313_D), .S(I_443_D));
  generic_nmos I_3440(.D(I_3440_D), .G(I_3441_G), .S(I_3440_S));
  generic_pmos I_3441(.D(I_3441_D), .G(I_3441_G), .S(I_3441_S));
  generic_nmos I_3442(.D(VSS), .G(I_3503_D), .S(I_3443_S));
  generic_pmos I_3443(.D(VDD), .G(I_3503_D), .S(I_3443_S));
  generic_nmos I_3444(.D(VSS), .G(I_3735_G), .S(I_3445_S));
  generic_pmos I_3445(.D(VDD), .G(I_3735_G), .S(I_3445_S));
  generic_nmos I_3446(.D(I_3446_D), .G(I_3511_S), .S(VSS));
  generic_pmos I_3447(.D(I_3447_D), .G(I_3511_S), .S(VDD));
  generic_nmos I_3448(.D(I_3448_D), .G(I_3607_D), .S(VSS));
  generic_pmos I_3449(.D(I_3449_D), .G(I_3607_D), .S(VDD));
  generic_pmos I_345(.D(VDD), .G(I_313_D), .S(I_443_D));
  generic_nmos I_3450(.D(I_3450_D), .G(I_3515_S), .S(VSS));
  generic_pmos I_3451(.D(I_3451_D), .G(I_3515_S), .S(VDD));
  generic_nmos I_3452(.D(I_3452_D), .G(I_3611_D), .S(VSS));
  generic_pmos I_3453(.D(I_3453_D), .G(I_3611_D), .S(VDD));
  generic_nmos I_3454(.D(VSS), .G(I_3455_G), .S(I_3454_S));
  generic_pmos I_3455(.D(VDD), .G(I_3455_G), .S(I_3455_S));
  generic_nmos I_3456(.D(I_3457_D), .G(I_3521_D), .S(I_3489_D));
  generic_pmos I_3457(.D(I_3457_D), .G(I_3555_G), .S(I_3489_D));
  generic_nmos I_3458(.D(VSS), .G(I_3427_D), .S(I_3491_S));
  generic_pmos I_3459(.D(VDD), .G(I_3587_D), .S(I_3491_D));
  generic_nmos I_346(.D(I_347_D), .G(I_603_D), .S(VSS));
  generic_nmos I_3460(.D(I_3461_D), .G(I_3333_S), .S(I_3493_D));
  generic_pmos I_3461(.D(I_3461_D), .G(I_3271_S), .S(I_3493_D));
  generic_nmos I_3462(.D(I_3493_S), .G(I_3271_S), .S(I_3495_D));
  generic_pmos I_3463(.D(I_3493_S), .G(I_3333_S), .S(I_3495_D));
  generic_nmos I_3464(.D(I_3591_S), .G(I_3499_D), .S(I_3497_S));
  generic_pmos I_3465(.D(I_3465_D), .G(I_3433_S), .S(I_3591_S));
  generic_nmos I_3466(.D(I_3499_D), .G(I_3497_S), .S(I_3499_S));
  generic_pmos I_3467(.D(I_3467_D), .G(I_3435_S), .S(I_3499_D));
  generic_nmos I_3468(.D(I_3501_D), .G(I_3597_S), .S(I_3500_D));
  generic_pmos I_3469(.D(VDD), .G(I_3431_S), .S(I_3501_D));
  generic_pmos I_347(.D(I_347_D), .G(I_603_D), .S(VDD));
  generic_nmos I_3470(.D(I_3471_D), .G(I_3407_D), .S(I_3503_D));
  generic_pmos I_3471(.D(I_3471_D), .G(I_3439_S), .S(I_3503_D));
  generic_nmos I_3472(.D(I_3505_D), .G(I_2319_D), .S(I_3504_D));
  generic_pmos I_3473(.D(VDD), .G(I_3663_S), .S(I_3505_D));
  generic_nmos I_3474(.D(I_3507_D), .G(I_3503_D), .S(I_3827_D));
  generic_pmos I_3475(.D(I_3475_D), .G(I_3443_S), .S(I_3507_D));
  generic_nmos I_3476(.D(I_3476_D), .G(I_3476_G), .S(I_3508_D));
  generic_pmos I_3477(.D(I_3477_D), .G(I_3508_G), .S(I_3509_D));
  generic_nmos I_3478(.D(I_3511_S), .G(I_3510_S), .S(VSS));
  generic_pmos I_3479(.D(I_3510_S), .G(I_1821_D), .S(VDD));
  generic_nmos I_348(.D(I_477_S), .G(I_317_D), .S(VSS));
  generic_nmos I_3480(.D(I_3480_D), .G(I_3480_G), .S(I_3512_D));
  generic_pmos I_3481(.D(I_3481_D), .G(I_3512_G), .S(I_3513_D));
  generic_nmos I_3482(.D(I_3515_S), .G(I_3514_S), .S(VSS));
  generic_pmos I_3483(.D(I_3514_S), .G(I_1821_D), .S(VDD));
  generic_nmos I_3484(.D(VSS), .G(I_3549_D), .S(I_3516_D));
  generic_pmos I_3485(.D(VDD), .G(I_3773_D), .S(I_3517_D));
  generic_nmos I_3486(.D(VSS), .G(I_3677_D), .S(I_3519_D));
  generic_pmos I_3487(.D(VDD), .G(I_3677_D), .S(I_3519_D));
  generic_nmos I_3488(.D(I_3489_D), .G(I_3555_G), .S(I_3489_S));
  generic_pmos I_3489(.D(I_3489_D), .G(I_3521_D), .S(I_3489_S));
  generic_pmos I_349(.D(I_477_S), .G(I_317_D), .S(VDD));
  generic_nmos I_3490(.D(I_3491_S), .G(I_3587_D), .S(VSS));
  generic_pmos I_3491(.D(I_3491_D), .G(I_3427_D), .S(I_3491_S));
  generic_nmos I_3492(.D(I_3493_D), .G(I_3271_S), .S(I_3493_S));
  generic_pmos I_3493(.D(I_3493_D), .G(I_3333_S), .S(I_3493_S));
  generic_nmos I_3494(.D(I_3495_D), .G(I_3333_S), .S(I_3495_S));
  generic_pmos I_3495(.D(I_3495_D), .G(I_3271_S), .S(I_3495_S));
  generic_nmos I_3496(.D(I_3497_S), .G(I_3433_S), .S(VSS));
  generic_pmos I_3497(.D(I_3591_S), .G(I_3433_S), .S(I_3497_S));
  generic_nmos I_3498(.D(I_3499_S), .G(I_3435_S), .S(VSS));
  generic_pmos I_3499(.D(I_3499_D), .G(I_3435_S), .S(I_3499_S));
  generic_pmos I_35(.D(VDD), .G(I_3_D), .S(I_67_D));
  generic_nmos I_350(.D(I_447_D), .G(I_319_D), .S(I_382_D));
  generic_nmos I_3500(.D(I_3500_D), .G(I_3431_S), .S(VSS));
  generic_pmos I_3501(.D(I_3501_D), .G(I_3597_S), .S(VDD));
  generic_nmos I_3502(.D(I_3503_D), .G(I_3439_S), .S(I_3503_S));
  generic_pmos I_3503(.D(I_3503_D), .G(I_3407_D), .S(I_3503_S));
  generic_nmos I_3504(.D(I_3504_D), .G(I_3663_S), .S(VSS));
  generic_pmos I_3505(.D(I_3505_D), .G(I_2319_D), .S(VDD));
  generic_nmos I_3506(.D(I_3827_D), .G(I_3443_S), .S(VSS));
  generic_pmos I_3507(.D(I_3507_D), .G(I_3443_S), .S(I_3827_D));
  generic_nmos I_3508(.D(I_3508_D), .G(I_3508_G), .S(I_3508_S));
  generic_pmos I_3509(.D(I_3509_D), .G(I_3509_G), .S(I_3509_S));
  generic_pmos I_351(.D(VDD), .G(I_319_D), .S(I_447_D));
  generic_nmos I_3510(.D(VSS), .G(I_1821_D), .S(I_3510_S));
  generic_pmos I_3511(.D(VDD), .G(I_3510_S), .S(I_3511_S));
  generic_nmos I_3512(.D(I_3512_D), .G(I_3512_G), .S(I_3512_S));
  generic_pmos I_3513(.D(I_3513_D), .G(I_3513_G), .S(I_3513_S));
  generic_nmos I_3514(.D(VSS), .G(I_1821_D), .S(I_3514_S));
  generic_pmos I_3515(.D(VDD), .G(I_3514_S), .S(I_3515_S));
  generic_nmos I_3516(.D(I_3516_D), .G(I_3773_D), .S(I_3517_D));
  generic_pmos I_3517(.D(I_3517_D), .G(I_3549_D), .S(VDD));
  generic_nmos I_3518(.D(I_3519_D), .G(I_3677_D), .S(VSS));
  generic_pmos I_3519(.D(I_3519_D), .G(I_3677_D), .S(VDD));
  generic_nmos I_352(.D(VSS), .G(I_448_D), .S(I_385_D));
  generic_nmos I_3520(.D(I_3521_D), .G(I_3555_G), .S(VSS));
  generic_pmos I_3521(.D(I_3521_D), .G(I_3555_G), .S(VDD));
  generic_nmos I_3522(.D(I_3587_D), .G(I_3333_S), .S(I_3554_D));
  generic_pmos I_3523(.D(I_3587_D), .G(I_3333_S), .S(VDD));
  generic_nmos I_3524(.D(I_3621_D), .G(I_3655_S), .S(VSS));
  generic_pmos I_3525(.D(I_3621_D), .G(I_3655_S), .S(VDD));
  generic_nmos I_3526(.D(I_3653_S), .G(I_3591_S), .S(I_3558_D));
  generic_pmos I_3527(.D(VDD), .G(I_3591_S), .S(I_3653_S));
  generic_nmos I_3528(.D(I_3529_D), .G(I_3529_G), .S(VSS));
  generic_pmos I_3529(.D(I_3529_D), .G(I_3529_G), .S(VDD));
  generic_pmos I_353(.D(VDD), .G(I_448_D), .S(I_385_D));
  generic_nmos I_3530(.D(VSS), .G(I_3431_S), .S(I_3562_D));
  generic_pmos I_3531(.D(I_3562_D), .G(I_3431_S), .S(I_3563_D));
  generic_nmos I_3532(.D(I_3565_D), .G(I_3499_S), .S(I_3564_D));
  generic_pmos I_3533(.D(VDD), .G(I_3499_S), .S(I_3565_D));
  generic_nmos I_3534(.D(I_3535_D), .G(I_3599_S), .S(VSS));
  generic_pmos I_3535(.D(I_3535_D), .G(I_3599_S), .S(VDD));
  generic_nmos I_3536(.D(VSS), .G(I_2319_D), .S(I_3568_D));
  generic_pmos I_3537(.D(I_3568_D), .G(I_2319_D), .S(I_3569_D));
  generic_nmos I_3538(.D(I_3538_D), .G(I_3539_G), .S(I_3570_D));
  generic_pmos I_3539(.D(I_3539_D), .G(I_3539_G), .S(I_3571_D));
  generic_nmos I_354(.D(I_354_D), .G(I_1249_D), .S(VSS));
  generic_nmos I_3540(.D(I_3540_D), .G(I_3541_G), .S(I_3572_D));
  generic_pmos I_3541(.D(I_3541_D), .G(I_3541_G), .S(I_3573_D));
  generic_nmos I_3542(.D(I_3607_D), .G(I_3351_S), .S(I_3574_D));
  generic_pmos I_3543(.D(I_3607_D), .G(I_3351_S), .S(VDD));
  generic_nmos I_3544(.D(I_3609_D), .G(I_3027_D), .S(I_3576_D));
  generic_pmos I_3545(.D(I_3609_D), .G(I_3027_D), .S(VDD));
  generic_nmos I_3546(.D(I_3611_D), .G(I_3355_S), .S(I_3578_D));
  generic_pmos I_3547(.D(I_3611_D), .G(I_3355_S), .S(VDD));
  generic_nmos I_3548(.D(I_3549_D), .G(I_1689_D), .S(VSS));
  generic_pmos I_3549(.D(I_3549_D), .G(I_1689_D), .S(VDD));
  generic_pmos I_355(.D(I_355_D), .G(I_1249_D), .S(VDD));
  generic_nmos I_3550(.D(I_3615_D), .G(I_3029_D), .S(I_3582_D));
  generic_pmos I_3551(.D(I_3615_D), .G(I_3029_D), .S(VDD));
  generic_nmos I_3552(.D(VSS), .G(I_3913_S), .S(I_3584_D));
  generic_pmos I_3553(.D(VDD), .G(I_3913_S), .S(I_3585_D));
  generic_nmos I_3554(.D(I_3554_D), .G(I_3555_G), .S(I_3586_D));
  generic_pmos I_3555(.D(VDD), .G(I_3555_G), .S(I_3587_D));
  generic_nmos I_3556(.D(VSS), .G(I_3241_D), .S(I_3588_D));
  generic_pmos I_3557(.D(VDD), .G(I_3241_D), .S(I_3655_S));
  generic_nmos I_3558(.D(I_3558_D), .G(I_3241_D), .S(VSS));
  generic_pmos I_3559(.D(I_3653_S), .G(I_3241_D), .S(VDD));
  generic_nmos I_356(.D(I_356_D), .G(I_389_S), .S(VSS));
  generic_nmos I_3560(.D(VSS), .G(I_3561_G), .S(VSS));
  generic_pmos I_3561(.D(VDD), .G(I_3561_G), .S(VDD));
  generic_nmos I_3562(.D(I_3562_D), .G(I_3657_D), .S(VSS));
  generic_pmos I_3563(.D(I_3563_D), .G(I_3657_D), .S(VDD));
  generic_nmos I_3564(.D(I_3564_D), .G(I_2253_D), .S(VSS));
  generic_pmos I_3565(.D(I_3565_D), .G(I_2253_D), .S(VDD));
  generic_nmos I_3566(.D(VSS), .G(I_3567_G), .S(VSS));
  generic_pmos I_3567(.D(VDD), .G(I_3567_G), .S(VDD));
  generic_nmos I_3568(.D(I_3568_D), .G(I_3663_S), .S(VSS));
  generic_pmos I_3569(.D(I_3569_D), .G(I_3663_S), .S(VDD));
  generic_pmos I_357(.D(I_421_D), .G(I_389_S), .S(VDD));
  generic_nmos I_3570(.D(I_3570_D), .G(I_3571_G), .S(I_3602_D));
  generic_pmos I_3571(.D(I_3571_D), .G(I_3571_G), .S(I_3603_D));
  generic_nmos I_3572(.D(I_3572_D), .G(I_3573_G), .S(I_3604_D));
  generic_pmos I_3573(.D(I_3573_D), .G(I_3573_G), .S(I_3605_D));
  generic_nmos I_3574(.D(I_3574_D), .G(I_3510_S), .S(I_3606_D));
  generic_pmos I_3575(.D(VDD), .G(I_3510_S), .S(I_3607_D));
  generic_nmos I_3576(.D(I_3576_D), .G(I_3832_S), .S(I_3608_D));
  generic_pmos I_3577(.D(VDD), .G(I_3832_S), .S(I_3609_D));
  generic_nmos I_3578(.D(I_3578_D), .G(I_3514_S), .S(I_3610_D));
  generic_pmos I_3579(.D(VDD), .G(I_3514_S), .S(I_3611_D));
  generic_nmos I_358(.D(VSS), .G(I_1187_S), .S(I_390_D));
  generic_nmos I_3580(.D(VSS), .G(I_1689_D), .S(I_3612_D));
  generic_pmos I_3581(.D(VDD), .G(I_1689_D), .S(I_3613_D));
  generic_nmos I_3582(.D(I_3582_D), .G(I_3838_S), .S(I_3614_D));
  generic_pmos I_3583(.D(VDD), .G(I_3838_S), .S(I_3615_D));
  generic_nmos I_3584(.D(I_3584_D), .G(I_3975_D), .S(I_3585_D));
  generic_pmos I_3585(.D(I_3585_D), .G(I_3975_D), .S(VDD));
  generic_nmos I_3586(.D(I_3586_D), .G(I_3173_S), .S(VSS));
  generic_pmos I_3587(.D(I_3587_D), .G(I_3173_S), .S(VDD));
  generic_nmos I_3588(.D(I_3588_D), .G(I_3653_D), .S(I_3655_S));
  generic_pmos I_3589(.D(I_3655_S), .G(I_3653_D), .S(VDD));
  generic_pmos I_359(.D(VDD), .G(I_1187_S), .S(I_453_S));
  generic_nmos I_3590(.D(VSS), .G(I_3655_D), .S(I_3591_S));
  generic_pmos I_3591(.D(VDD), .G(I_3655_D), .S(I_3591_S));
  generic_nmos I_3592(.D(VSS), .G(I_3593_G), .S(I_3593_S));
  generic_pmos I_3593(.D(VDD), .G(I_3593_G), .S(I_3593_S));
  generic_nmos I_3594(.D(VSS), .G(I_3593_S), .S(I_3595_S));
  generic_pmos I_3595(.D(VDD), .G(I_3593_S), .S(I_3595_S));
  generic_nmos I_3596(.D(VSS), .G(I_2253_D), .S(I_3597_S));
  generic_pmos I_3597(.D(VDD), .G(I_2253_D), .S(I_3597_S));
  generic_nmos I_3598(.D(VSS), .G(I_3825_D), .S(I_3599_S));
  generic_pmos I_3599(.D(VDD), .G(I_3825_D), .S(I_3599_S));
  generic_nmos I_36(.D(I_36_D), .G(I_69_S), .S(VSS));
  generic_nmos I_360(.D(VSS), .G(I_361_G), .S(VSS));
  generic_nmos I_3600(.D(VSS), .G(I_3568_D), .S(I_3601_S));
  generic_pmos I_3601(.D(VDD), .G(I_3568_D), .S(I_3601_S));
  generic_nmos I_3602(.D(I_3602_D), .G(I_3603_G), .S(I_3602_S));
  generic_pmos I_3603(.D(I_3603_D), .G(I_3603_G), .S(I_3603_S));
  generic_nmos I_3604(.D(I_3604_D), .G(I_3605_G), .S(I_3604_S));
  generic_pmos I_3605(.D(I_3605_D), .G(I_3605_G), .S(I_3605_S));
  generic_nmos I_3606(.D(I_3606_D), .G(I_1962_D), .S(VSS));
  generic_pmos I_3607(.D(I_3607_D), .G(I_1962_D), .S(VDD));
  generic_nmos I_3608(.D(I_3608_D), .G(I_3672_S), .S(VSS));
  generic_pmos I_3609(.D(I_3609_D), .G(I_3672_S), .S(VDD));
  generic_pmos I_361(.D(VDD), .G(I_361_G), .S(VDD));
  generic_nmos I_3610(.D(I_3610_D), .G(VDD), .S(VSS));
  generic_pmos I_3611(.D(I_3611_D), .G(VDD), .S(VDD));
  generic_nmos I_3612(.D(I_3612_D), .G(I_3997_D), .S(I_3613_D));
  generic_pmos I_3613(.D(I_3613_D), .G(I_3997_D), .S(VDD));
  generic_nmos I_3614(.D(I_3614_D), .G(I_3678_S), .S(VSS));
  generic_pmos I_3615(.D(I_3615_D), .G(I_3678_S), .S(VDD));
  generic_nmos I_3616(.D(VSS), .G(I_3649_G), .S(I_3649_D));
  generic_pmos I_3617(.D(VDD), .G(I_3649_G), .S(I_3649_D));
  generic_nmos I_3618(.D(VSS), .G(I_3755_S), .S(I_3651_D));
  generic_pmos I_3619(.D(VDD), .G(I_3755_S), .S(I_3651_D));
  generic_nmos I_362(.D(I_362_D), .G(I_297_S), .S(I_394_D));
  generic_nmos I_3620(.D(I_3621_D), .G(I_3493_S), .S(I_3653_D));
  generic_pmos I_3621(.D(I_3621_D), .G(I_3431_S), .S(I_3653_D));
  generic_nmos I_3622(.D(I_3653_S), .G(I_3431_S), .S(I_3655_D));
  generic_pmos I_3623(.D(I_3653_S), .G(I_3493_S), .S(I_3655_D));
  generic_nmos I_3624(.D(VSS), .G(I_3813_S), .S(I_3657_D));
  generic_pmos I_3625(.D(VDD), .G(I_3813_S), .S(I_3657_D));
  generic_nmos I_3626(.D(I_3659_S), .G(I_3659_G), .S(VSS));
  generic_pmos I_3627(.D(I_3627_D), .G(I_3658_G), .S(VDD));
  generic_nmos I_3628(.D(I_3725_D), .G(I_3595_S), .S(I_3660_D));
  generic_pmos I_3629(.D(I_3725_D), .G(I_3919_S), .S(VDD));
  generic_pmos I_363(.D(VDD), .G(I_297_S), .S(I_395_D));
  generic_nmos I_3630(.D(I_3759_S), .G(I_3823_D), .S(I_3663_D));
  generic_pmos I_3631(.D(I_3759_S), .G(I_3695_D), .S(I_3663_D));
  generic_nmos I_3632(.D(VSS), .G(I_3568_D), .S(I_3825_D));
  generic_pmos I_3633(.D(I_3633_D), .G(I_3664_G), .S(I_3825_D));
  generic_nmos I_3634(.D(I_3763_S), .G(I_3827_D), .S(I_3667_D));
  generic_pmos I_3635(.D(I_3763_S), .G(I_3699_D), .S(I_3667_D));
  generic_nmos I_3636(.D(I_3765_S), .G(I_3829_D), .S(I_3669_D));
  generic_pmos I_3637(.D(I_3765_S), .G(I_3701_D), .S(I_3669_D));
  generic_nmos I_3638(.D(I_3638_D), .G(I_3638_G), .S(I_3670_D));
  generic_pmos I_3639(.D(I_3639_D), .G(I_3670_G), .S(I_3671_D));
  generic_nmos I_364(.D(I_364_D), .G(I_365_G), .S(I_396_D));
  generic_nmos I_3640(.D(I_3673_S), .G(I_3672_S), .S(VSS));
  generic_pmos I_3641(.D(I_3672_S), .G(I_1597_D), .S(VDD));
  generic_nmos I_3642(.D(VSS), .G(I_3995_D), .S(I_3675_D));
  generic_pmos I_3643(.D(VDD), .G(I_3995_D), .S(I_3675_D));
  generic_nmos I_3644(.D(I_3677_D), .G(I_3613_D), .S(I_3676_D));
  generic_pmos I_3645(.D(VDD), .G(I_3517_D), .S(I_3677_D));
  generic_nmos I_3646(.D(I_3679_S), .G(I_3678_S), .S(VSS));
  generic_pmos I_3647(.D(I_3678_S), .G(I_1597_D), .S(VDD));
  generic_nmos I_3648(.D(I_3649_D), .G(I_3649_G), .S(VSS));
  generic_pmos I_3649(.D(I_3649_D), .G(I_3649_G), .S(VDD));
  generic_pmos I_365(.D(I_365_D), .G(I_365_G), .S(I_397_D));
  generic_nmos I_3650(.D(I_3651_D), .G(I_3755_S), .S(VSS));
  generic_pmos I_3651(.D(I_3651_D), .G(I_3755_S), .S(VDD));
  generic_nmos I_3652(.D(I_3653_D), .G(I_3431_S), .S(I_3653_S));
  generic_pmos I_3653(.D(I_3653_D), .G(I_3493_S), .S(I_3653_S));
  generic_nmos I_3654(.D(I_3655_D), .G(I_3493_S), .S(I_3655_S));
  generic_pmos I_3655(.D(I_3655_D), .G(I_3431_S), .S(I_3655_S));
  generic_nmos I_3656(.D(I_3657_D), .G(I_3813_S), .S(VSS));
  generic_pmos I_3657(.D(I_3657_D), .G(I_3813_S), .S(VDD));
  generic_nmos I_3658(.D(VSS), .G(I_3658_G), .S(I_3658_S));
  generic_pmos I_3659(.D(VDD), .G(I_3659_G), .S(I_3659_S));
  generic_nmos I_366(.D(I_366_D), .G(I_367_G), .S(I_398_D));
  generic_nmos I_3660(.D(I_3660_D), .G(I_3919_S), .S(I_3692_D));
  generic_pmos I_3661(.D(VDD), .G(I_3595_S), .S(I_3725_D));
  generic_nmos I_3662(.D(I_3663_D), .G(I_3695_D), .S(I_3663_S));
  generic_pmos I_3663(.D(I_3663_D), .G(I_3823_D), .S(I_3663_S));
  generic_nmos I_3664(.D(I_3825_D), .G(I_3664_G), .S(I_3664_S));
  generic_pmos I_3665(.D(I_3825_D), .G(I_3505_D), .S(VDD));
  generic_nmos I_3666(.D(I_3667_D), .G(I_3699_D), .S(I_3667_S));
  generic_pmos I_3667(.D(I_3667_D), .G(I_3827_D), .S(I_3667_S));
  generic_nmos I_3668(.D(I_3669_D), .G(I_3701_D), .S(I_3669_S));
  generic_pmos I_3669(.D(I_3669_D), .G(I_3829_D), .S(I_3669_S));
  generic_pmos I_367(.D(I_367_D), .G(I_367_G), .S(I_399_D));
  generic_nmos I_3670(.D(I_3670_D), .G(I_3670_G), .S(I_3670_S));
  generic_pmos I_3671(.D(I_3671_D), .G(I_3671_G), .S(I_3671_S));
  generic_nmos I_3672(.D(VSS), .G(I_1597_D), .S(I_3672_S));
  generic_pmos I_3673(.D(VDD), .G(I_3672_S), .S(I_3673_S));
  generic_nmos I_3674(.D(I_3675_D), .G(I_3995_D), .S(VSS));
  generic_pmos I_3675(.D(I_3675_D), .G(I_3995_D), .S(VDD));
  generic_nmos I_3676(.D(I_3676_D), .G(I_3517_D), .S(VSS));
  generic_pmos I_3677(.D(I_3677_D), .G(I_3613_D), .S(VDD));
  generic_nmos I_3678(.D(VSS), .G(I_1597_D), .S(I_3678_S));
  generic_pmos I_3679(.D(VDD), .G(I_3678_S), .S(I_3679_S));
  generic_nmos I_368(.D(I_368_D), .G(I_369_G), .S(I_400_D));
  generic_nmos I_3680(.D(I_3681_D), .G(I_3649_D), .S(VSS));
  generic_pmos I_3681(.D(I_3681_D), .G(I_3649_D), .S(VDD));
  generic_nmos I_3682(.D(I_3683_D), .G(I_3649_D), .S(VSS));
  generic_pmos I_3683(.D(I_3683_D), .G(I_3649_D), .S(VDD));
  generic_nmos I_3684(.D(I_3781_D), .G(I_3815_S), .S(VSS));
  generic_pmos I_3685(.D(I_3781_D), .G(I_3815_S), .S(VDD));
  generic_nmos I_3686(.D(I_3813_S), .G(I_3751_S), .S(I_3718_D));
  generic_pmos I_3687(.D(VDD), .G(I_3751_S), .S(I_3813_S));
  generic_nmos I_3688(.D(I_3753_D), .G(I_3915_G), .S(I_3720_D));
  generic_pmos I_3689(.D(I_3753_D), .G(I_3915_G), .S(VDD));
  generic_pmos I_369(.D(I_369_D), .G(I_369_G), .S(I_401_D));
  generic_nmos I_3690(.D(I_3691_D), .G(I_3659_S), .S(VSS));
  generic_pmos I_3691(.D(I_3691_D), .G(I_3659_S), .S(VDD));
  generic_nmos I_3692(.D(I_3692_D), .G(I_3691_D), .S(I_3724_D));
  generic_pmos I_3693(.D(VDD), .G(I_3691_D), .S(I_3725_D));
  generic_nmos I_3694(.D(I_3695_D), .G(I_3823_D), .S(VSS));
  generic_pmos I_3695(.D(I_3695_D), .G(I_3823_D), .S(VDD));
  generic_nmos I_3696(.D(I_3985_S), .G(I_3601_S), .S(I_3728_D));
  generic_pmos I_3697(.D(VDD), .G(I_3601_S), .S(I_3985_S));
  generic_nmos I_3698(.D(I_3699_D), .G(I_3827_D), .S(VSS));
  generic_pmos I_3699(.D(I_3699_D), .G(I_3827_D), .S(VDD));
  generic_pmos I_37(.D(I_101_D), .G(I_69_S), .S(VDD));
  generic_nmos I_370(.D(I_370_D), .G(I_371_G), .S(I_402_D));
  generic_nmos I_3700(.D(I_3701_D), .G(I_3829_D), .S(VSS));
  generic_pmos I_3701(.D(I_3701_D), .G(I_3829_D), .S(VDD));
  generic_nmos I_3702(.D(I_3703_D), .G(I_3735_G), .S(VSS));
  generic_pmos I_3703(.D(I_3703_D), .G(I_3735_G), .S(VDD));
  generic_nmos I_3704(.D(I_3769_D), .G(I_3990_S), .S(I_3736_D));
  generic_pmos I_3705(.D(I_3769_D), .G(I_3990_S), .S(VDD));
  generic_nmos I_3706(.D(I_3771_D), .G(I_3609_D), .S(I_3738_D));
  generic_pmos I_3707(.D(I_3771_D), .G(I_3609_D), .S(VDD));
  generic_nmos I_3708(.D(I_3773_D), .G(I_3615_D), .S(I_3740_D));
  generic_pmos I_3709(.D(I_3773_D), .G(I_3615_D), .S(VDD));
  generic_pmos I_371(.D(I_371_D), .G(I_371_G), .S(I_403_D));
  generic_nmos I_3710(.D(I_3775_D), .G(I_3988_S), .S(I_3742_D));
  generic_pmos I_3711(.D(I_3775_D), .G(I_3988_S), .S(VDD));
  generic_nmos I_3712(.D(VSS), .G(I_3649_D), .S(I_3744_D));
  generic_pmos I_3713(.D(VDD), .G(I_3649_D), .S(I_3745_D));
  generic_nmos I_3714(.D(VSS), .G(I_3649_D), .S(I_3746_D));
  generic_pmos I_3715(.D(VDD), .G(I_3649_D), .S(I_3747_D));
  generic_nmos I_3716(.D(VSS), .G(I_3241_D), .S(I_3748_D));
  generic_pmos I_3717(.D(VDD), .G(I_3241_D), .S(I_3815_S));
  generic_nmos I_3718(.D(I_3718_D), .G(I_3241_D), .S(VSS));
  generic_pmos I_3719(.D(I_3813_S), .G(I_3241_D), .S(VDD));
  generic_nmos I_372(.D(I_372_D), .G(I_437_D), .S(VSS));
  generic_nmos I_3720(.D(I_3720_D), .G(I_3969_S), .S(I_3752_D));
  generic_pmos I_3721(.D(VDD), .G(I_3969_S), .S(I_3753_D));
  generic_nmos I_3722(.D(VSS), .G(I_3725_D), .S(I_3755_S));
  generic_pmos I_3723(.D(VDD), .G(I_3725_D), .S(I_3755_D));
  generic_nmos I_3724(.D(I_3724_D), .G(I_3859_D), .S(VSS));
  generic_pmos I_3725(.D(I_3725_D), .G(I_3859_D), .S(VDD));
  generic_nmos I_3726(.D(VSS), .G(I_3727_G), .S(VSS));
  generic_pmos I_3727(.D(VDD), .G(I_3727_G), .S(VDD));
  generic_nmos I_3728(.D(I_3728_D), .G(I_3505_D), .S(VSS));
  generic_pmos I_3729(.D(I_3985_S), .G(I_3505_D), .S(VDD));
  generic_pmos I_373(.D(I_373_D), .G(I_437_D), .S(VDD));
  generic_nmos I_3730(.D(VSS), .G(I_3731_G), .S(VSS));
  generic_pmos I_3731(.D(VDD), .G(I_3731_G), .S(VDD));
  generic_nmos I_3732(.D(VSS), .G(I_3733_G), .S(VSS));
  generic_pmos I_3733(.D(VDD), .G(I_3733_G), .S(VDD));
  generic_nmos I_3734(.D(VSS), .G(I_3735_G), .S(I_3766_D));
  generic_pmos I_3735(.D(VDD), .G(I_3735_G), .S(I_3767_D));
  generic_nmos I_3736(.D(I_3736_D), .G(I_3672_S), .S(I_3768_D));
  generic_pmos I_3737(.D(VDD), .G(I_3672_S), .S(I_3769_D));
  generic_nmos I_3738(.D(I_3738_D), .G(I_3769_D), .S(I_3770_D));
  generic_pmos I_3739(.D(VDD), .G(I_3769_D), .S(I_3771_D));
  generic_nmos I_374(.D(I_375_D), .G(I_471_D), .S(VSS));
  generic_nmos I_3740(.D(I_3740_D), .G(I_3775_D), .S(I_3772_D));
  generic_pmos I_3741(.D(VDD), .G(I_3775_D), .S(I_3773_D));
  generic_nmos I_3742(.D(I_3742_D), .G(I_3678_S), .S(I_3774_D));
  generic_pmos I_3743(.D(VDD), .G(I_3678_S), .S(I_3775_D));
  generic_nmos I_3744(.D(I_3744_D), .G(I_2791_S), .S(I_3745_D));
  generic_pmos I_3745(.D(I_3745_D), .G(I_2791_S), .S(VDD));
  generic_nmos I_3746(.D(I_3746_D), .G(I_1741_S), .S(I_3747_D));
  generic_pmos I_3747(.D(I_3747_D), .G(I_1741_S), .S(VDD));
  generic_nmos I_3748(.D(I_3748_D), .G(I_3813_D), .S(I_3815_S));
  generic_pmos I_3749(.D(I_3815_S), .G(I_3813_D), .S(VDD));
  generic_pmos I_375(.D(I_375_D), .G(I_471_D), .S(VDD));
  generic_nmos I_3750(.D(VSS), .G(I_3815_D), .S(I_3751_S));
  generic_pmos I_3751(.D(VDD), .G(I_3815_D), .S(I_3751_S));
  generic_nmos I_3752(.D(I_3752_D), .G(I_3847_G), .S(VSS));
  generic_pmos I_3753(.D(I_3753_D), .G(I_3847_G), .S(VDD));
  generic_nmos I_3754(.D(I_3755_S), .G(I_3883_D), .S(VSS));
  generic_pmos I_3755(.D(I_3755_D), .G(I_3883_D), .S(I_3755_S));
  generic_nmos I_3756(.D(VSS), .G(I_3659_S), .S(I_3788_D));
  generic_pmos I_3757(.D(VDD), .G(I_3659_S), .S(I_3884_D));
  generic_nmos I_3758(.D(VSS), .G(I_3663_S), .S(I_3759_S));
  generic_pmos I_3759(.D(VDD), .G(I_3663_S), .S(I_3759_S));
  generic_nmos I_376(.D(I_443_D), .G(I_313_D), .S(VSS));
  generic_nmos I_3760(.D(VSS), .G(I_3985_S), .S(I_3953_D));
  generic_pmos I_3761(.D(VDD), .G(I_3985_S), .S(I_3953_D));
  generic_nmos I_3762(.D(VSS), .G(I_3667_S), .S(I_3763_S));
  generic_pmos I_3763(.D(VDD), .G(I_3667_S), .S(I_3763_S));
  generic_nmos I_3764(.D(VSS), .G(I_3669_S), .S(I_3765_S));
  generic_pmos I_3765(.D(VDD), .G(I_3669_S), .S(I_3765_S));
  generic_nmos I_3766(.D(I_3766_D), .G(I_3767_G), .S(I_3767_D));
  generic_pmos I_3767(.D(I_3767_D), .G(I_3767_G), .S(VDD));
  generic_nmos I_3768(.D(I_3768_D), .G(I_3833_S), .S(VSS));
  generic_pmos I_3769(.D(I_3769_D), .G(I_3833_S), .S(VDD));
  generic_pmos I_377(.D(I_443_D), .G(I_313_D), .S(VDD));
  generic_nmos I_3770(.D(I_3770_D), .G(I_3929_D), .S(VSS));
  generic_pmos I_3771(.D(I_3771_D), .G(I_3929_D), .S(VDD));
  generic_nmos I_3772(.D(I_3772_D), .G(I_3935_D), .S(VSS));
  generic_pmos I_3773(.D(I_3773_D), .G(I_3935_D), .S(VDD));
  generic_nmos I_3774(.D(I_3774_D), .G(I_3839_S), .S(VSS));
  generic_pmos I_3775(.D(I_3775_D), .G(I_3839_S), .S(VDD));
  generic_nmos I_3776(.D(VSS), .G(I_3681_D), .S(I_3808_D));
  generic_pmos I_3777(.D(VDD), .G(I_2631_S), .S(I_3809_D));
  generic_nmos I_3778(.D(VSS), .G(I_3683_D), .S(I_3810_D));
  generic_pmos I_3779(.D(VDD), .G(I_2791_S), .S(I_3811_D));
  generic_nmos I_378(.D(VSS), .G(I_379_G), .S(I_410_D));
  generic_nmos I_3780(.D(I_3781_D), .G(I_3653_S), .S(I_3813_D));
  generic_pmos I_3781(.D(I_3781_D), .G(I_3591_S), .S(I_3813_D));
  generic_nmos I_3782(.D(I_3813_S), .G(I_3591_S), .S(I_3815_D));
  generic_pmos I_3783(.D(I_3813_S), .G(I_3653_S), .S(I_3815_D));
  generic_nmos I_3784(.D(I_3817_D), .G(I_3847_D), .S(I_3816_D));
  generic_pmos I_3785(.D(VDD), .G(I_3977_G), .S(I_3817_D));
  generic_nmos I_3786(.D(I_3883_D), .G(I_3819_G), .S(I_3818_D));
  generic_pmos I_3787(.D(I_3883_D), .G(I_3988_S), .S(VDD));
  generic_nmos I_3788(.D(I_3788_D), .G(I_3983_D), .S(I_3820_D));
  generic_pmos I_3789(.D(VDD), .G(I_3977_G), .S(I_3884_D));
  generic_pmos I_379(.D(VDD), .G(I_379_G), .S(I_411_D));
  generic_nmos I_3790(.D(I_3823_D), .G(I_3663_S), .S(I_3823_S));
  generic_pmos I_3791(.D(I_3791_D), .G(I_3759_S), .S(I_3823_D));
  generic_nmos I_3792(.D(I_3825_D), .G(I_3953_D), .S(I_3825_S));
  generic_pmos I_3793(.D(I_3793_D), .G(I_3824_G), .S(I_3825_D));
  generic_nmos I_3794(.D(I_3827_D), .G(I_3667_S), .S(I_3829_D));
  generic_pmos I_3795(.D(I_3795_D), .G(I_3763_S), .S(I_3827_D));
  generic_nmos I_3796(.D(I_3829_D), .G(I_3669_S), .S(I_3829_S));
  generic_pmos I_3797(.D(I_3797_D), .G(I_3765_S), .S(I_3829_D));
  generic_nmos I_3798(.D(VSS), .G(I_3703_D), .S(I_3830_D));
  generic_pmos I_3799(.D(VDD), .G(I_3830_G), .S(I_3831_D));
  generic_nmos I_38(.D(VSS), .G(I_1187_S), .S(I_70_D));
  generic_nmos I_380(.D(VSS), .G(I_381_G), .S(VSS));
  generic_nmos I_3800(.D(I_3833_S), .G(I_3832_S), .S(VSS));
  generic_pmos I_3801(.D(I_3832_S), .G(I_1821_D), .S(VDD));
  generic_nmos I_3802(.D(VSS), .G(I_3867_D), .S(I_3834_D));
  generic_pmos I_3803(.D(VDD), .G(I_3771_D), .S(I_3835_D));
  generic_nmos I_3804(.D(VSS), .G(I_3869_D), .S(I_3836_D));
  generic_pmos I_3805(.D(VDD), .G(I_3836_G), .S(I_3837_D));
  generic_nmos I_3806(.D(I_3839_S), .G(I_3838_S), .S(VSS));
  generic_pmos I_3807(.D(I_3838_S), .G(I_1821_D), .S(VDD));
  generic_nmos I_3808(.D(I_3808_D), .G(I_2631_S), .S(I_3809_D));
  generic_pmos I_3809(.D(I_3809_D), .G(I_3681_D), .S(VDD));
  generic_pmos I_381(.D(VDD), .G(I_381_G), .S(VDD));
  generic_nmos I_3810(.D(I_3810_D), .G(I_2791_S), .S(I_3811_D));
  generic_pmos I_3811(.D(I_3811_D), .G(I_3683_D), .S(VDD));
  generic_nmos I_3812(.D(I_3813_D), .G(I_3591_S), .S(I_3813_S));
  generic_pmos I_3813(.D(I_3813_D), .G(I_3653_S), .S(I_3813_S));
  generic_nmos I_3814(.D(I_3815_D), .G(I_3653_S), .S(I_3815_S));
  generic_pmos I_3815(.D(I_3815_D), .G(I_3591_S), .S(I_3815_S));
  generic_nmos I_3816(.D(I_3816_D), .G(I_3977_G), .S(VSS));
  generic_pmos I_3817(.D(I_3817_D), .G(I_3847_D), .S(VDD));
  generic_nmos I_3818(.D(I_3818_D), .G(I_3988_S), .S(I_3850_D));
  generic_pmos I_3819(.D(VDD), .G(I_3819_G), .S(I_3883_D));
  generic_nmos I_382(.D(I_382_D), .G(I_639_S), .S(VSS));
  generic_nmos I_3820(.D(I_3820_D), .G(I_3977_G), .S(I_3852_D));
  generic_pmos I_3821(.D(I_3884_D), .G(I_3983_D), .S(VDD));
  generic_nmos I_3822(.D(I_3823_S), .G(I_3759_S), .S(VSS));
  generic_pmos I_3823(.D(I_3823_D), .G(I_3759_S), .S(I_3823_S));
  generic_nmos I_3824(.D(I_3825_S), .G(I_3824_G), .S(I_3824_S));
  generic_pmos I_3825(.D(I_3825_D), .G(I_3985_S), .S(I_3825_S));
  generic_nmos I_3826(.D(I_3829_D), .G(I_3763_S), .S(VSS));
  generic_pmos I_3827(.D(I_3827_D), .G(I_3763_S), .S(I_3829_D));
  generic_nmos I_3828(.D(I_3829_S), .G(I_3765_S), .S(VSS));
  generic_pmos I_3829(.D(I_3829_D), .G(I_3765_S), .S(I_3829_S));
  generic_pmos I_383(.D(I_447_D), .G(I_639_S), .S(VDD));
  generic_nmos I_3830(.D(I_3830_D), .G(I_3830_G), .S(I_3831_D));
  generic_pmos I_3831(.D(I_3831_D), .G(I_3703_D), .S(VDD));
  generic_nmos I_3832(.D(VSS), .G(I_1821_D), .S(I_3832_S));
  generic_pmos I_3833(.D(VDD), .G(I_3832_S), .S(I_3833_S));
  generic_nmos I_3834(.D(I_3834_D), .G(I_3771_D), .S(I_3835_D));
  generic_pmos I_3835(.D(I_3835_D), .G(I_3867_D), .S(VDD));
  generic_nmos I_3836(.D(I_3836_D), .G(I_3836_G), .S(I_3837_D));
  generic_pmos I_3837(.D(I_3837_D), .G(I_3869_D), .S(VDD));
  generic_nmos I_3838(.D(VSS), .G(I_1821_D), .S(I_3838_S));
  generic_pmos I_3839(.D(VDD), .G(I_3838_S), .S(I_3839_S));
  generic_nmos I_384(.D(I_385_D), .G(I_448_D), .S(VSS));
  generic_nmos I_3840(.D(VSS), .G(I_3745_D), .S(I_3872_D));
  generic_pmos I_3841(.D(VDD), .G(I_3745_D), .S(I_3904_D));
  generic_nmos I_3842(.D(VSS), .G(I_3747_D), .S(I_3874_D));
  generic_pmos I_3843(.D(VDD), .G(I_3747_D), .S(I_3906_D));
  generic_nmos I_3844(.D(I_3845_D), .G(I_3649_D), .S(VSS));
  generic_pmos I_3845(.D(I_3845_D), .G(I_3649_D), .S(VDD));
  generic_nmos I_3846(.D(I_3847_D), .G(I_3847_G), .S(VSS));
  generic_pmos I_3847(.D(I_3847_D), .G(I_3847_G), .S(VDD));
  generic_nmos I_3848(.D(VSS), .G(I_3817_D), .S(I_3880_D));
  generic_pmos I_3849(.D(VDD), .G(I_3817_D), .S(I_3913_S));
  generic_pmos I_385(.D(I_385_D), .G(I_448_D), .S(VDD));
  generic_nmos I_3850(.D(I_3850_D), .G(I_3851_G), .S(I_3882_D));
  generic_pmos I_3851(.D(VDD), .G(I_3851_G), .S(I_3883_D));
  generic_nmos I_3852(.D(I_3852_D), .G(I_3529_D), .S(I_3884_D));
  generic_pmos I_3853(.D(I_3884_D), .G(I_3529_D), .S(VDD));
  generic_nmos I_3854(.D(I_3854_D), .G(I_3855_G), .S(I_3887_D));
  generic_pmos I_3855(.D(I_3855_D), .G(I_3855_G), .S(I_3887_D));
  generic_nmos I_3856(.D(I_3856_D), .G(I_3857_G), .S(I_3889_D));
  generic_pmos I_3857(.D(I_3857_D), .G(I_3857_G), .S(I_3889_D));
  generic_nmos I_3858(.D(I_3859_D), .G(I_3923_S), .S(VSS));
  generic_pmos I_3859(.D(I_3859_D), .G(I_3923_S), .S(VDD));
  generic_nmos I_386(.D(VSS), .G(I_1249_D), .S(I_387_S));
  generic_nmos I_3860(.D(I_3861_D), .G(I_3195_S), .S(VSS));
  generic_pmos I_3861(.D(I_3861_D), .G(I_3195_S), .S(VDD));
  generic_nmos I_3862(.D(VSS), .G(I_3767_D), .S(I_3894_D));
  generic_pmos I_3863(.D(VDD), .G(I_3767_D), .S(I_3926_D));
  generic_nmos I_3864(.D(I_3929_D), .G(I_3673_S), .S(I_3896_D));
  generic_pmos I_3865(.D(I_3929_D), .G(I_3673_S), .S(VDD));
  generic_nmos I_3866(.D(I_3867_D), .G(I_1689_D), .S(VSS));
  generic_pmos I_3867(.D(I_3867_D), .G(I_1689_D), .S(VDD));
  generic_nmos I_3868(.D(I_3869_D), .G(I_1755_D), .S(VSS));
  generic_pmos I_3869(.D(I_3869_D), .G(I_1755_D), .S(VDD));
  generic_pmos I_387(.D(VDD), .G(I_1249_D), .S(I_387_S));
  generic_nmos I_3870(.D(I_3935_D), .G(I_3679_S), .S(I_3902_D));
  generic_pmos I_3871(.D(I_3935_D), .G(I_3679_S), .S(VDD));
  generic_nmos I_3872(.D(I_3872_D), .G(I_3809_D), .S(I_3904_D));
  generic_pmos I_3873(.D(I_3904_D), .G(I_3809_D), .S(VDD));
  generic_nmos I_3874(.D(I_3874_D), .G(I_3811_D), .S(I_3906_D));
  generic_pmos I_3875(.D(I_3906_D), .G(I_3811_D), .S(VDD));
  generic_nmos I_3876(.D(VSS), .G(I_3649_D), .S(I_3908_D));
  generic_pmos I_3877(.D(VDD), .G(I_3649_D), .S(I_3909_D));
  generic_nmos I_3878(.D(VSS), .G(I_3845_D), .S(I_3910_D));
  generic_pmos I_3879(.D(VDD), .G(I_3845_D), .S(I_3911_D));
  generic_nmos I_388(.D(VSS), .G(I_453_D), .S(I_389_S));
  generic_nmos I_3880(.D(I_3880_D), .G(I_3753_D), .S(I_3912_D));
  generic_pmos I_3881(.D(I_3913_S), .G(I_3753_D), .S(VDD));
  generic_nmos I_3882(.D(I_3882_D), .G(I_3887_D), .S(VSS));
  generic_pmos I_3883(.D(I_3883_D), .G(I_3887_D), .S(VDD));
  generic_nmos I_3884(.D(I_3884_D), .G(VSS), .S(VSS));
  generic_pmos I_3885(.D(VDD), .G(VSS), .S(VDD));
  generic_nmos I_3886(.D(I_3887_D), .G(I_3987_S), .S(VSS));
  generic_pmos I_3887(.D(I_3887_D), .G(I_3987_S), .S(VDD));
  generic_nmos I_3888(.D(I_3889_D), .G(I_3825_S), .S(VSS));
  generic_pmos I_3889(.D(I_3889_D), .G(I_3825_S), .S(VDD));
  generic_pmos I_389(.D(VDD), .G(I_453_D), .S(I_389_S));
  generic_nmos I_3890(.D(VSS), .G(I_3861_D), .S(VSS));
  generic_pmos I_3891(.D(VDD), .G(I_3861_D), .S(VDD));
  generic_nmos I_3892(.D(VSS), .G(I_3893_G), .S(I_3924_D));
  generic_pmos I_3893(.D(VDD), .G(I_3893_G), .S(I_3925_D));
  generic_nmos I_3894(.D(I_3894_D), .G(I_3831_D), .S(I_3926_D));
  generic_pmos I_3895(.D(I_3926_D), .G(I_3831_D), .S(VDD));
  generic_nmos I_3896(.D(I_3896_D), .G(I_3832_S), .S(I_3928_D));
  generic_pmos I_3897(.D(VDD), .G(I_3832_S), .S(I_3929_D));
  generic_nmos I_3898(.D(VSS), .G(I_1689_D), .S(I_3930_D));
  generic_pmos I_3899(.D(VDD), .G(I_1689_D), .S(I_3931_D));
  generic_pmos I_39(.D(VDD), .G(I_1187_S), .S(I_133_S));
  generic_nmos I_390(.D(I_390_D), .G(I_455_D), .S(I_453_S));
  generic_nmos I_3900(.D(VSS), .G(I_1755_D), .S(I_3932_D));
  generic_pmos I_3901(.D(VDD), .G(I_1755_D), .S(I_3933_D));
  generic_nmos I_3902(.D(I_3902_D), .G(I_3838_S), .S(I_3934_D));
  generic_pmos I_3903(.D(VDD), .G(I_3838_S), .S(I_3935_D));
  generic_nmos I_3904(.D(I_3904_D), .G(I_3905_G), .S(I_3904_S));
  generic_pmos I_3905(.D(VDD), .G(I_3905_G), .S(I_3905_S));
  generic_nmos I_3906(.D(I_3906_D), .G(I_3907_G), .S(I_3906_S));
  generic_pmos I_3907(.D(VDD), .G(I_3907_G), .S(I_3907_S));
  generic_nmos I_3908(.D(I_3908_D), .G(I_2631_S), .S(I_3909_D));
  generic_pmos I_3909(.D(I_3909_D), .G(I_2631_S), .S(VDD));
  generic_pmos I_391(.D(I_453_S), .G(I_455_D), .S(VDD));
  generic_nmos I_3910(.D(I_3910_D), .G(I_3911_G), .S(I_3911_D));
  generic_pmos I_3911(.D(I_3911_D), .G(I_3911_G), .S(VDD));
  generic_nmos I_3912(.D(I_3912_D), .G(I_3977_D), .S(I_3913_S));
  generic_pmos I_3913(.D(VDD), .G(I_3977_D), .S(I_3913_S));
  generic_nmos I_3914(.D(VSS), .G(I_3915_G), .S(I_3915_S));
  generic_pmos I_3915(.D(VDD), .G(I_3915_G), .S(I_3915_S));
  generic_nmos I_3916(.D(VSS), .G(I_3529_D), .S(I_3917_S));
  generic_pmos I_3917(.D(VDD), .G(I_3529_D), .S(I_3917_S));
  generic_nmos I_3918(.D(VSS), .G(I_3983_D), .S(I_3919_S));
  generic_pmos I_3919(.D(VDD), .G(I_3983_D), .S(I_3919_S));
  generic_nmos I_392(.D(VSS), .G(I_555_D), .S(I_393_S));
  generic_nmos I_3920(.D(VSS), .G(I_3889_D), .S(I_3921_S));
  generic_pmos I_3921(.D(VDD), .G(I_3889_D), .S(I_3921_S));
  generic_nmos I_3922(.D(VSS), .G(I_3923_G), .S(I_3923_S));
  generic_pmos I_3923(.D(VDD), .G(I_3923_G), .S(I_3923_S));
  generic_nmos I_3924(.D(I_3924_D), .G(I_3925_G), .S(I_3924_S));
  generic_pmos I_3925(.D(I_3925_D), .G(I_3925_G), .S(I_3925_S));
  generic_nmos I_3926(.D(I_3926_D), .G(I_3927_G), .S(I_3926_S));
  generic_pmos I_3927(.D(VDD), .G(I_3927_G), .S(I_3927_S));
  generic_nmos I_3928(.D(I_3928_D), .G(I_3129_D), .S(VSS));
  generic_pmos I_3929(.D(I_3929_D), .G(I_3129_D), .S(VDD));
  generic_pmos I_393(.D(VDD), .G(I_555_D), .S(I_393_S));
  generic_nmos I_3930(.D(I_3930_D), .G(I_3926_D), .S(I_3931_D));
  generic_pmos I_3931(.D(I_3931_D), .G(I_3926_D), .S(VDD));
  generic_nmos I_3932(.D(I_3932_D), .G(I_3933_G), .S(I_3933_D));
  generic_pmos I_3933(.D(I_3933_D), .G(I_3933_G), .S(VDD));
  generic_nmos I_3934(.D(I_3934_D), .G(I_2969_D), .S(VSS));
  generic_pmos I_3935(.D(I_3935_D), .G(I_2969_D), .S(VDD));
  generic_nmos I_3936(.D(I_3969_S), .G(I_3971_S), .S(VSS));
  generic_pmos I_3937(.D(I_3937_D), .G(I_3968_G), .S(VDD));
  generic_nmos I_3938(.D(I_3971_S), .G(I_3971_G), .S(VSS));
  generic_pmos I_3939(.D(I_3939_D), .G(I_3970_G), .S(VDD));
  generic_nmos I_394(.D(I_394_D), .G(I_461_S), .S(VSS));
  generic_nmos I_3940(.D(I_3973_D), .G(I_3909_D), .S(I_3972_D));
  generic_pmos I_3941(.D(VDD), .G(I_3911_D), .S(I_3973_D));
  generic_nmos I_3942(.D(VSS), .G(I_3755_S), .S(I_3974_D));
  generic_pmos I_3943(.D(VDD), .G(I_3974_G), .S(I_3975_D));
  generic_nmos I_3944(.D(I_3977_D), .G(I_3977_G), .S(I_3976_D));
  generic_pmos I_3945(.D(VDD), .G(I_3915_S), .S(I_3977_D));
  generic_nmos I_3946(.D(VSS), .G(I_3981_D), .S(I_3979_D));
  generic_pmos I_3947(.D(VDD), .G(I_3981_D), .S(I_3979_D));
  generic_nmos I_3948(.D(I_3981_D), .G(I_3917_S), .S(I_3980_D));
  generic_pmos I_3949(.D(VDD), .G(I_3980_G), .S(I_3981_D));
  generic_pmos I_395(.D(I_395_D), .G(I_461_S), .S(VDD));
  generic_nmos I_3950(.D(I_3950_D), .G(I_3950_G), .S(VSS));
  generic_pmos I_3951(.D(VDD), .G(I_3982_G), .S(I_3983_D));
  generic_nmos I_3952(.D(I_3953_D), .G(I_3889_D), .S(I_3985_D));
  generic_pmos I_3953(.D(I_3953_D), .G(I_3921_S), .S(I_3985_D));
  generic_nmos I_3954(.D(I_3987_S), .G(I_3987_G), .S(VSS));
  generic_pmos I_3955(.D(I_3955_D), .G(I_3986_G), .S(VDD));
  generic_nmos I_3956(.D(I_3956_D), .G(I_3956_G), .S(VSS));
  generic_pmos I_3957(.D(I_3988_S), .G(I_3988_G), .S(VDD));
  generic_nmos I_3958(.D(I_3958_D), .G(I_3958_G), .S(VSS));
  generic_pmos I_3959(.D(I_3990_S), .G(I_3990_G), .S(VDD));
  generic_nmos I_396(.D(I_396_D), .G(I_397_G), .S(I_396_S));
  generic_nmos I_3960(.D(I_3993_S), .G(I_3993_G), .S(VSS));
  generic_pmos I_3961(.D(I_3961_D), .G(I_3992_G), .S(VDD));
  generic_nmos I_3962(.D(I_3995_D), .G(I_3931_D), .S(I_3994_D));
  generic_pmos I_3963(.D(VDD), .G(I_3835_D), .S(I_3995_D));
  generic_nmos I_3964(.D(I_3997_D), .G(I_3933_D), .S(I_3996_D));
  generic_pmos I_3965(.D(VDD), .G(I_3837_D), .S(I_3997_D));
  generic_nmos I_3966(.D(VSS), .G(I_3999_G), .S(I_3999_D));
  generic_pmos I_3967(.D(VDD), .G(I_3999_G), .S(I_3999_D));
  generic_nmos I_3968(.D(VSS), .G(I_3968_G), .S(I_3968_S));
  generic_pmos I_3969(.D(VDD), .G(I_3971_S), .S(I_3969_S));
  generic_pmos I_397(.D(I_397_D), .G(I_397_G), .S(I_397_S));
  generic_nmos I_3970(.D(VSS), .G(I_3970_G), .S(I_3970_S));
  generic_pmos I_3971(.D(VDD), .G(I_3971_G), .S(I_3971_S));
  generic_nmos I_3972(.D(I_3972_D), .G(I_3911_D), .S(VSS));
  generic_pmos I_3973(.D(I_3973_D), .G(I_3909_D), .S(VDD));
  generic_nmos I_3974(.D(I_3974_D), .G(I_3974_G), .S(I_3975_D));
  generic_pmos I_3975(.D(I_3975_D), .G(I_3755_S), .S(VDD));
  generic_nmos I_3976(.D(I_3976_D), .G(I_3915_S), .S(VSS));
  generic_pmos I_3977(.D(I_3977_D), .G(I_3977_G), .S(VDD));
  generic_nmos I_3978(.D(I_3979_D), .G(I_3981_D), .S(VSS));
  generic_pmos I_3979(.D(I_3979_D), .G(I_3981_D), .S(VDD));
  generic_nmos I_398(.D(I_398_D), .G(I_399_G), .S(I_398_S));
  generic_nmos I_3980(.D(I_3980_D), .G(I_3980_G), .S(VSS));
  generic_pmos I_3981(.D(I_3981_D), .G(I_3917_S), .S(VDD));
  generic_nmos I_3982(.D(VSS), .G(I_3982_G), .S(I_3983_D));
  generic_pmos I_3983(.D(I_3983_D), .G(I_3983_G), .S(I_3983_S));
  generic_nmos I_3984(.D(I_3985_D), .G(I_3921_S), .S(I_3985_S));
  generic_pmos I_3985(.D(I_3985_D), .G(I_3889_D), .S(I_3985_S));
  generic_nmos I_3986(.D(VSS), .G(I_3986_G), .S(I_3986_S));
  generic_pmos I_3987(.D(VDD), .G(I_3987_G), .S(I_3987_S));
  generic_nmos I_3988(.D(VSS), .G(I_3988_G), .S(I_3988_S));
  generic_pmos I_3989(.D(VDD), .G(I_3989_G), .S(I_3989_S));
  generic_pmos I_399(.D(I_399_D), .G(I_399_G), .S(I_399_S));
  generic_nmos I_3990(.D(VSS), .G(I_3990_G), .S(I_3990_S));
  generic_pmos I_3991(.D(VDD), .G(I_3991_G), .S(I_3991_S));
  generic_nmos I_3992(.D(VSS), .G(I_3992_G), .S(I_3992_S));
  generic_pmos I_3993(.D(VDD), .G(I_3993_G), .S(I_3993_S));
  generic_nmos I_3994(.D(I_3994_D), .G(I_3835_D), .S(VSS));
  generic_pmos I_3995(.D(I_3995_D), .G(I_3931_D), .S(VDD));
  generic_nmos I_3996(.D(I_3996_D), .G(I_3837_D), .S(VSS));
  generic_pmos I_3997(.D(I_3997_D), .G(I_3933_D), .S(VDD));
  generic_nmos I_3998(.D(I_3999_D), .G(I_3999_G), .S(VSS));
  generic_pmos I_3999(.D(I_3999_D), .G(I_3999_G), .S(VDD));
  generic_nmos I_4(.D(I_101_D), .G(I_1187_S), .S(I_36_D));
  generic_nmos I_40(.D(I_40_D), .G(I_41_G), .S(I_72_D));
  generic_nmos I_400(.D(I_400_D), .G(I_401_G), .S(I_400_S));
  generic_pmos I_401(.D(I_401_D), .G(I_401_G), .S(I_401_S));
  generic_nmos I_402(.D(I_402_D), .G(I_403_G), .S(I_402_S));
  generic_pmos I_403(.D(I_403_D), .G(I_403_G), .S(I_403_S));
  generic_nmos I_404(.D(VSS), .G(I_405_G), .S(I_404_S));
  generic_pmos I_405(.D(VDD), .G(I_405_G), .S(I_405_S));
  generic_nmos I_406(.D(VSS), .G(I_375_D), .S(I_439_D));
  generic_pmos I_407(.D(VDD), .G(I_375_D), .S(I_439_D));
  generic_nmos I_408(.D(VSS), .G(I_443_D), .S(I_409_S));
  generic_pmos I_409(.D(VDD), .G(I_443_D), .S(I_409_S));
  generic_pmos I_41(.D(I_41_D), .G(I_41_G), .S(I_73_D));
  generic_nmos I_410(.D(I_410_D), .G(I_411_G), .S(I_410_S));
  generic_pmos I_411(.D(I_411_D), .G(I_411_G), .S(I_411_S));
  generic_nmos I_412(.D(VSS), .G(I_477_S), .S(I_445_D));
  generic_pmos I_413(.D(VDD), .G(I_477_S), .S(I_445_D));
  generic_nmos I_414(.D(VSS), .G(I_447_D), .S(I_415_S));
  generic_pmos I_415(.D(VDD), .G(I_447_D), .S(I_415_S));
  generic_nmos I_416(.D(VSS), .G(I_545_D), .S(I_448_D));
  generic_pmos I_417(.D(I_448_D), .G(I_1089_D), .S(I_449_D));
  generic_nmos I_418(.D(I_418_D), .G(I_418_G), .S(I_450_D));
  generic_pmos I_419(.D(I_419_D), .G(I_450_G), .S(I_451_D));
  generic_nmos I_42(.D(I_42_D), .G(I_43_G), .S(I_74_D));
  generic_nmos I_420(.D(I_421_D), .G(I_329_D), .S(I_453_D));
  generic_pmos I_421(.D(I_421_D), .G(I_395_D), .S(I_453_D));
  generic_nmos I_422(.D(I_423_D), .G(I_395_D), .S(I_455_D));
  generic_pmos I_423(.D(I_423_D), .G(I_329_D), .S(I_455_D));
  generic_nmos I_424(.D(I_457_D), .G(I_2905_D), .S(I_456_D));
  generic_pmos I_425(.D(VDD), .G(I_3065_D), .S(I_457_D));
  generic_nmos I_426(.D(I_426_D), .G(I_426_G), .S(VSS));
  generic_pmos I_427(.D(I_458_S), .G(I_461_S), .S(VDD));
  generic_nmos I_428(.D(I_461_S), .G(I_2809_D), .S(VSS));
  generic_pmos I_429(.D(I_429_D), .G(I_460_G), .S(VDD));
  generic_pmos I_43(.D(I_43_D), .G(I_43_G), .S(I_75_D));
  generic_nmos I_430(.D(I_430_D), .G(I_430_G), .S(I_462_D));
  generic_pmos I_431(.D(I_431_D), .G(I_462_G), .S(I_463_D));
  generic_nmos I_432(.D(I_432_D), .G(I_432_G), .S(I_464_D));
  generic_pmos I_433(.D(I_433_D), .G(I_464_G), .S(I_465_D));
  generic_nmos I_434(.D(I_434_D), .G(I_434_G), .S(I_466_D));
  generic_pmos I_435(.D(I_435_D), .G(I_466_G), .S(I_467_D));
  generic_nmos I_436(.D(I_437_D), .G(I_1373_S), .S(I_468_D));
  generic_pmos I_437(.D(I_437_D), .G(I_1373_S), .S(I_469_D));
  generic_nmos I_438(.D(I_439_D), .G(I_251_S), .S(I_471_D));
  generic_pmos I_439(.D(I_439_D), .G(I_315_D), .S(I_471_D));
  generic_nmos I_44(.D(I_44_D), .G(I_45_G), .S(I_76_D));
  generic_nmos I_440(.D(I_475_D), .G(I_315_D), .S(I_473_D));
  generic_pmos I_441(.D(I_475_D), .G(I_251_S), .S(I_473_D));
  generic_nmos I_442(.D(I_443_D), .G(I_789_D), .S(I_475_D));
  generic_pmos I_443(.D(I_443_D), .G(I_1045_D), .S(I_475_D));
  generic_nmos I_444(.D(I_445_D), .G(I_509_D), .S(I_477_D));
  generic_pmos I_445(.D(I_445_D), .G(I_573_D), .S(I_477_D));
  generic_nmos I_446(.D(I_447_D), .G(I_95_D), .S(I_479_D));
  generic_pmos I_447(.D(I_447_D), .G(I_93_S), .S(I_479_D));
  generic_nmos I_448(.D(I_448_D), .G(I_1089_D), .S(VSS));
  generic_pmos I_449(.D(I_449_D), .G(I_545_D), .S(VDD));
  generic_pmos I_45(.D(I_45_D), .G(I_45_G), .S(I_77_D));
  generic_nmos I_450(.D(I_450_D), .G(I_450_G), .S(I_450_S));
  generic_pmos I_451(.D(I_451_D), .G(I_451_G), .S(I_451_S));
  generic_nmos I_452(.D(I_453_D), .G(I_395_D), .S(I_453_S));
  generic_pmos I_453(.D(I_453_D), .G(I_329_D), .S(I_453_S));
  generic_nmos I_454(.D(I_455_D), .G(I_329_D), .S(I_1415_S));
  generic_pmos I_455(.D(I_455_D), .G(I_395_D), .S(I_1415_S));
  generic_nmos I_456(.D(I_456_D), .G(I_3065_D), .S(VSS));
  generic_pmos I_457(.D(I_457_D), .G(I_2905_D), .S(VDD));
  generic_nmos I_458(.D(VSS), .G(I_461_S), .S(I_458_S));
  generic_pmos I_459(.D(VDD), .G(I_459_G), .S(I_459_S));
  generic_nmos I_46(.D(I_46_D), .G(I_47_G), .S(I_78_D));
  generic_nmos I_460(.D(VSS), .G(I_460_G), .S(I_460_S));
  generic_pmos I_461(.D(VDD), .G(I_2809_D), .S(I_461_S));
  generic_nmos I_462(.D(I_462_D), .G(I_462_G), .S(I_462_S));
  generic_pmos I_463(.D(I_463_D), .G(I_463_G), .S(I_463_S));
  generic_nmos I_464(.D(I_464_D), .G(I_464_G), .S(I_464_S));
  generic_pmos I_465(.D(I_465_D), .G(I_465_G), .S(I_465_S));
  generic_nmos I_466(.D(I_466_D), .G(I_466_G), .S(I_466_S));
  generic_pmos I_467(.D(I_467_D), .G(I_467_G), .S(I_467_S));
  generic_nmos I_468(.D(I_468_D), .G(I_1373_S), .S(VSS));
  generic_pmos I_469(.D(I_469_D), .G(I_1373_S), .S(VDD));
  generic_pmos I_47(.D(I_47_D), .G(I_47_G), .S(I_79_D));
  generic_nmos I_470(.D(I_471_D), .G(I_315_D), .S(I_471_S));
  generic_pmos I_471(.D(I_471_D), .G(I_251_S), .S(I_471_S));
  generic_nmos I_472(.D(I_473_D), .G(I_251_S), .S(I_505_D));
  generic_pmos I_473(.D(I_473_D), .G(I_315_D), .S(I_505_D));
  generic_nmos I_474(.D(I_475_D), .G(I_1045_D), .S(I_2201_D));
  generic_pmos I_475(.D(I_475_D), .G(I_789_D), .S(I_2201_D));
  generic_nmos I_476(.D(I_477_D), .G(I_573_D), .S(I_477_S));
  generic_pmos I_477(.D(I_477_D), .G(I_509_D), .S(I_477_S));
  generic_nmos I_478(.D(I_479_D), .G(I_93_S), .S(I_575_S));
  generic_pmos I_479(.D(I_479_D), .G(I_95_D), .S(I_575_S));
  generic_nmos I_48(.D(I_48_D), .G(I_49_G), .S(I_80_D));
  generic_nmos I_480(.D(I_544_D), .G(I_1832_D), .S(I_545_D));
  generic_pmos I_481(.D(VDD), .G(I_1832_D), .S(I_513_D));
  generic_nmos I_482(.D(I_482_D), .G(I_483_G), .S(VSS));
  generic_pmos I_483(.D(I_483_D), .G(I_483_G), .S(VDD));
  generic_nmos I_484(.D(I_581_D), .G(I_1187_S), .S(I_516_D));
  generic_pmos I_485(.D(VDD), .G(I_1187_S), .S(I_581_D));
  generic_nmos I_486(.D(I_583_D), .G(I_613_S), .S(VSS));
  generic_pmos I_487(.D(I_583_D), .G(I_613_S), .S(VDD));
  generic_nmos I_488(.D(I_553_D), .G(I_524_D), .S(I_520_D));
  generic_pmos I_489(.D(I_553_D), .G(I_524_D), .S(VDD));
  generic_pmos I_49(.D(I_49_D), .G(I_49_G), .S(I_81_D));
  generic_nmos I_490(.D(I_555_D), .G(I_458_S), .S(I_522_D));
  generic_pmos I_491(.D(I_555_D), .G(I_458_S), .S(VDD));
  generic_nmos I_492(.D(VSS), .G(I_493_G), .S(I_524_D));
  generic_pmos I_493(.D(I_524_D), .G(I_493_G), .S(I_525_D));
  generic_nmos I_494(.D(I_494_D), .G(I_495_G), .S(I_526_D));
  generic_pmos I_495(.D(I_495_D), .G(I_495_G), .S(I_527_D));
  generic_nmos I_496(.D(I_496_D), .G(I_497_G), .S(I_528_D));
  generic_pmos I_497(.D(I_497_D), .G(I_497_G), .S(I_529_D));
  generic_nmos I_498(.D(I_498_D), .G(I_499_G), .S(I_530_D));
  generic_pmos I_499(.D(I_499_D), .G(I_499_G), .S(I_531_D));
  generic_pmos I_5(.D(VDD), .G(I_1187_S), .S(I_101_D));
  generic_nmos I_50(.D(I_50_D), .G(I_51_G), .S(I_82_D));
  generic_nmos I_500(.D(I_500_D), .G(I_501_G), .S(I_532_D));
  generic_pmos I_501(.D(I_501_D), .G(I_501_G), .S(I_533_D));
  generic_nmos I_502(.D(I_503_D), .G(I_503_G), .S(VSS));
  generic_pmos I_503(.D(I_503_D), .G(I_503_G), .S(VDD));
  generic_nmos I_504(.D(I_505_D), .G(I_601_D), .S(VSS));
  generic_pmos I_505(.D(I_505_D), .G(I_601_D), .S(VDD));
  generic_nmos I_506(.D(I_2201_D), .G(I_507_G), .S(VSS));
  generic_pmos I_507(.D(I_2201_D), .G(I_507_G), .S(VDD));
  generic_nmos I_508(.D(I_509_D), .G(I_573_D), .S(VSS));
  generic_pmos I_509(.D(I_509_D), .G(I_573_D), .S(VDD));
  generic_pmos I_51(.D(I_51_D), .G(I_51_G), .S(I_83_D));
  generic_nmos I_510(.D(I_511_D), .G(I_479_D), .S(VSS));
  generic_pmos I_511(.D(I_511_D), .G(I_479_D), .S(VDD));
  generic_nmos I_512(.D(I_545_D), .G(I_547_D), .S(I_544_D));
  generic_pmos I_513(.D(I_513_D), .G(I_547_D), .S(I_545_D));
  generic_nmos I_514(.D(VSS), .G(I_611_D), .S(I_546_D));
  generic_pmos I_515(.D(VDD), .G(I_611_D), .S(I_547_D));
  generic_nmos I_516(.D(I_516_D), .G(I_549_S), .S(VSS));
  generic_pmos I_517(.D(I_581_D), .G(I_549_S), .S(VDD));
  generic_nmos I_518(.D(VSS), .G(I_1187_S), .S(I_550_D));
  generic_pmos I_519(.D(VDD), .G(I_1187_S), .S(I_613_S));
  generic_nmos I_52(.D(I_52_D), .G(I_53_G), .S(VSS));
  generic_nmos I_520(.D(I_520_D), .G(I_3065_D), .S(I_552_D));
  generic_pmos I_521(.D(VDD), .G(I_3065_D), .S(I_553_D));
  generic_nmos I_522(.D(I_522_D), .G(I_616_S), .S(I_554_D));
  generic_pmos I_523(.D(VDD), .G(I_616_S), .S(I_555_D));
  generic_nmos I_524(.D(I_524_D), .G(I_1211_D), .S(VSS));
  generic_pmos I_525(.D(I_525_D), .G(I_1211_D), .S(VDD));
  generic_nmos I_526(.D(I_526_D), .G(I_527_G), .S(I_558_D));
  generic_pmos I_527(.D(I_527_D), .G(I_527_G), .S(I_559_D));
  generic_nmos I_528(.D(I_528_D), .G(I_529_G), .S(I_560_D));
  generic_pmos I_529(.D(I_529_D), .G(I_529_G), .S(I_561_D));
  generic_pmos I_53(.D(I_53_D), .G(I_53_G), .S(VDD));
  generic_nmos I_530(.D(I_530_D), .G(I_531_G), .S(I_562_D));
  generic_pmos I_531(.D(I_531_D), .G(I_531_G), .S(I_563_D));
  generic_nmos I_532(.D(I_532_D), .G(I_533_G), .S(I_564_D));
  generic_pmos I_533(.D(I_533_D), .G(I_533_G), .S(I_565_D));
  generic_nmos I_534(.D(VSS), .G(I_535_G), .S(I_566_D));
  generic_pmos I_535(.D(VDD), .G(I_535_G), .S(I_567_D));
  generic_nmos I_536(.D(VSS), .G(I_473_D), .S(I_601_D));
  generic_pmos I_537(.D(VDD), .G(I_473_D), .S(I_601_D));
  generic_nmos I_538(.D(VSS), .G(I_539_G), .S(VSS));
  generic_pmos I_539(.D(VDD), .G(I_539_G), .S(VDD));
  generic_nmos I_54(.D(VSS), .G(I_55_G), .S(VSS));
  generic_nmos I_540(.D(VSS), .G(I_511_D), .S(I_572_D));
  generic_pmos I_541(.D(VDD), .G(I_511_D), .S(I_573_D));
  generic_nmos I_542(.D(VSS), .G(I_543_G), .S(VSS));
  generic_pmos I_543(.D(VDD), .G(I_543_G), .S(VDD));
  generic_nmos I_544(.D(I_544_D), .G(I_609_D), .S(VSS));
  generic_pmos I_545(.D(I_545_D), .G(I_609_D), .S(VDD));
  generic_nmos I_546(.D(I_546_D), .G(I_675_D), .S(I_547_D));
  generic_pmos I_547(.D(I_547_D), .G(I_675_D), .S(VDD));
  generic_nmos I_548(.D(VSS), .G(I_613_D), .S(I_549_S));
  generic_pmos I_549(.D(VDD), .G(I_613_D), .S(I_549_S));
  generic_pmos I_55(.D(VDD), .G(I_55_G), .S(VDD));
  generic_nmos I_550(.D(I_550_D), .G(I_615_D), .S(I_613_S));
  generic_pmos I_551(.D(I_613_S), .G(I_615_D), .S(VDD));
  generic_nmos I_552(.D(I_552_D), .G(I_2905_D), .S(VSS));
  generic_pmos I_553(.D(I_553_D), .G(I_2905_D), .S(VDD));
  generic_nmos I_554(.D(I_554_D), .G(I_618_S), .S(VSS));
  generic_pmos I_555(.D(I_555_D), .G(I_618_S), .S(VDD));
  generic_nmos I_556(.D(VSS), .G(I_557_G), .S(I_556_S));
  generic_pmos I_557(.D(VDD), .G(I_557_G), .S(I_557_S));
  generic_nmos I_558(.D(I_558_D), .G(I_559_G), .S(I_558_S));
  generic_pmos I_559(.D(I_559_D), .G(I_559_G), .S(I_559_S));
  generic_nmos I_56(.D(I_56_D), .G(I_57_G), .S(I_88_D));
  generic_nmos I_560(.D(I_560_D), .G(I_561_G), .S(I_560_S));
  generic_pmos I_561(.D(I_561_D), .G(I_561_G), .S(I_561_S));
  generic_nmos I_562(.D(I_562_D), .G(I_563_G), .S(I_562_S));
  generic_pmos I_563(.D(I_563_D), .G(I_563_G), .S(I_563_S));
  generic_nmos I_564(.D(I_564_D), .G(I_565_G), .S(I_564_S));
  generic_pmos I_565(.D(I_565_D), .G(I_565_G), .S(I_565_S));
  generic_nmos I_566(.D(I_566_D), .G(I_567_G), .S(I_566_S));
  generic_pmos I_567(.D(I_567_D), .G(I_567_G), .S(I_567_S));
  generic_nmos I_568(.D(I_601_D), .G(I_473_D), .S(VSS));
  generic_pmos I_569(.D(I_601_D), .G(I_473_D), .S(VDD));
  generic_pmos I_57(.D(I_57_D), .G(I_57_G), .S(I_89_D));
  generic_nmos I_570(.D(VSS), .G(I_571_G), .S(I_2841_D));
  generic_pmos I_571(.D(VDD), .G(I_571_G), .S(I_2841_D));
  generic_nmos I_572(.D(I_572_D), .G(I_957_S), .S(I_573_D));
  generic_pmos I_573(.D(I_573_D), .G(I_957_S), .S(VDD));
  generic_nmos I_574(.D(VSS), .G(I_511_D), .S(I_575_S));
  generic_pmos I_575(.D(VDD), .G(I_511_D), .S(I_575_S));
  generic_nmos I_576(.D(VSS), .G(I_547_D), .S(I_608_D));
  generic_pmos I_577(.D(VDD), .G(I_1832_D), .S(I_609_D));
  generic_nmos I_578(.D(I_611_D), .G(I_707_S), .S(I_610_D));
  generic_pmos I_579(.D(VDD), .G(I_709_S), .S(I_611_D));
  generic_nmos I_58(.D(I_59_D), .G(I_1115_D), .S(VSS));
  generic_nmos I_580(.D(I_581_D), .G(I_393_S), .S(I_613_D));
  generic_pmos I_581(.D(I_581_D), .G(I_555_D), .S(I_613_D));
  generic_nmos I_582(.D(I_583_D), .G(I_555_D), .S(I_615_D));
  generic_pmos I_583(.D(I_583_D), .G(I_393_S), .S(I_615_D));
  generic_nmos I_584(.D(I_584_D), .G(I_584_G), .S(VSS));
  generic_pmos I_585(.D(I_616_S), .G(I_2649_D), .S(VDD));
  generic_nmos I_586(.D(I_586_D), .G(I_586_G), .S(VSS));
  generic_pmos I_587(.D(I_618_S), .G(I_553_D), .S(VDD));
  generic_nmos I_588(.D(I_588_D), .G(I_588_G), .S(I_620_D));
  generic_pmos I_589(.D(I_589_D), .G(I_620_G), .S(I_621_D));
  generic_pmos I_59(.D(I_59_D), .G(I_1115_D), .S(VDD));
  generic_nmos I_590(.D(I_590_D), .G(I_590_G), .S(I_622_D));
  generic_pmos I_591(.D(I_591_D), .G(I_622_G), .S(I_623_D));
  generic_nmos I_592(.D(I_592_D), .G(I_592_G), .S(I_624_D));
  generic_pmos I_593(.D(I_593_D), .G(I_624_G), .S(I_625_D));
  generic_nmos I_594(.D(I_594_D), .G(I_594_G), .S(I_626_D));
  generic_pmos I_595(.D(I_595_D), .G(I_626_G), .S(I_627_D));
  generic_nmos I_596(.D(I_596_D), .G(I_596_G), .S(I_628_D));
  generic_pmos I_597(.D(I_597_D), .G(I_628_G), .S(I_629_D));
  generic_nmos I_598(.D(I_2841_D), .G(I_1045_D), .S(I_631_D));
  generic_pmos I_599(.D(I_2841_D), .G(I_789_D), .S(I_631_D));
  generic_nmos I_6(.D(I_103_D), .G(I_133_S), .S(VSS));
  generic_nmos I_60(.D(I_93_S), .G(I_503_G), .S(VSS));
  generic_nmos I_600(.D(I_601_D), .G(I_251_S), .S(I_633_D));
  generic_pmos I_601(.D(I_601_D), .G(I_315_D), .S(I_633_D));
  generic_nmos I_602(.D(I_603_D), .G(I_667_D), .S(I_634_D));
  generic_pmos I_603(.D(I_603_D), .G(I_667_D), .S(I_635_D));
  generic_nmos I_604(.D(I_957_D), .G(I_93_S), .S(I_637_D));
  generic_pmos I_605(.D(I_957_D), .G(I_95_D), .S(I_637_D));
  generic_nmos I_606(.D(I_1407_D), .G(I_93_S), .S(I_639_S));
  generic_pmos I_607(.D(I_607_D), .G(I_638_G), .S(I_1407_D));
  generic_nmos I_608(.D(I_608_D), .G(I_1832_D), .S(I_609_D));
  generic_pmos I_609(.D(I_609_D), .G(I_547_D), .S(VDD));
  generic_pmos I_61(.D(I_93_S), .G(I_503_G), .S(VDD));
  generic_nmos I_610(.D(I_610_D), .G(I_709_S), .S(VSS));
  generic_pmos I_611(.D(I_611_D), .G(I_707_S), .S(VDD));
  generic_nmos I_612(.D(I_613_D), .G(I_555_D), .S(I_613_S));
  generic_pmos I_613(.D(I_613_D), .G(I_393_S), .S(I_613_S));
  generic_nmos I_614(.D(I_615_D), .G(I_393_S), .S(I_2169_D));
  generic_pmos I_615(.D(I_615_D), .G(I_555_D), .S(I_2169_D));
  generic_nmos I_616(.D(VSS), .G(I_2649_D), .S(I_616_S));
  generic_pmos I_617(.D(VDD), .G(I_617_G), .S(I_617_S));
  generic_nmos I_618(.D(VSS), .G(I_553_D), .S(I_618_S));
  generic_pmos I_619(.D(VDD), .G(I_619_G), .S(I_619_S));
  generic_nmos I_62(.D(VSS), .G(I_95_G), .S(I_95_D));
  generic_nmos I_620(.D(I_620_D), .G(I_620_G), .S(I_620_S));
  generic_pmos I_621(.D(I_621_D), .G(I_621_G), .S(I_621_S));
  generic_nmos I_622(.D(I_622_D), .G(I_622_G), .S(I_622_S));
  generic_pmos I_623(.D(I_623_D), .G(I_623_G), .S(I_623_S));
  generic_nmos I_624(.D(I_624_D), .G(I_624_G), .S(I_624_S));
  generic_pmos I_625(.D(I_625_D), .G(I_625_G), .S(I_625_S));
  generic_nmos I_626(.D(I_626_D), .G(I_626_G), .S(I_626_S));
  generic_pmos I_627(.D(I_627_D), .G(I_627_G), .S(I_627_S));
  generic_nmos I_628(.D(I_628_D), .G(I_628_G), .S(I_628_S));
  generic_pmos I_629(.D(I_629_D), .G(I_629_G), .S(I_629_S));
  generic_pmos I_63(.D(VDD), .G(I_95_G), .S(I_95_D));
  generic_nmos I_630(.D(I_631_D), .G(I_789_D), .S(I_727_D));
  generic_pmos I_631(.D(I_631_D), .G(I_1045_D), .S(I_727_D));
  generic_nmos I_632(.D(I_633_D), .G(I_315_D), .S(I_729_S));
  generic_pmos I_633(.D(I_633_D), .G(I_251_S), .S(I_729_S));
  generic_nmos I_634(.D(I_634_D), .G(I_667_D), .S(VSS));
  generic_pmos I_635(.D(I_635_D), .G(I_667_D), .S(VDD));
  generic_nmos I_636(.D(I_637_D), .G(I_95_D), .S(I_733_S));
  generic_pmos I_637(.D(I_637_D), .G(I_93_S), .S(I_733_S));
  generic_nmos I_638(.D(I_639_S), .G(I_638_G), .S(I_638_S));
  generic_pmos I_639(.D(I_1407_D), .G(I_95_D), .S(I_639_S));
  generic_nmos I_64(.D(VSS), .G(I_128_D), .S(I_65_S));
  generic_nmos I_640(.D(I_640_D), .G(I_641_G), .S(VSS));
  generic_pmos I_641(.D(I_641_D), .G(I_641_G), .S(VDD));
  generic_nmos I_642(.D(I_675_D), .G(I_1189_D), .S(I_674_D));
  generic_pmos I_643(.D(VDD), .G(I_1189_D), .S(I_675_D));
  generic_nmos I_644(.D(I_741_D), .G(I_1187_S), .S(I_676_D));
  generic_pmos I_645(.D(VDD), .G(I_1187_S), .S(I_741_D));
  generic_nmos I_646(.D(I_743_D), .G(I_773_S), .S(VSS));
  generic_pmos I_647(.D(I_743_D), .G(I_773_S), .S(VDD));
  generic_nmos I_648(.D(I_648_D), .G(I_649_G), .S(I_680_D));
  generic_pmos I_649(.D(I_649_D), .G(I_649_G), .S(I_681_D));
  generic_pmos I_65(.D(VDD), .G(I_128_D), .S(I_65_S));
  generic_nmos I_650(.D(I_715_D), .G(I_461_S), .S(I_682_D));
  generic_pmos I_651(.D(I_715_D), .G(I_461_S), .S(VDD));
  generic_nmos I_652(.D(I_652_D), .G(I_653_G), .S(I_684_D));
  generic_pmos I_653(.D(I_653_D), .G(I_653_G), .S(I_685_D));
  generic_nmos I_654(.D(I_654_D), .G(I_655_G), .S(I_686_D));
  generic_pmos I_655(.D(I_655_D), .G(I_655_G), .S(I_687_D));
  generic_nmos I_656(.D(I_656_D), .G(I_657_G), .S(I_688_D));
  generic_pmos I_657(.D(I_657_D), .G(I_657_G), .S(I_689_D));
  generic_nmos I_658(.D(I_658_D), .G(I_659_G), .S(I_690_D));
  generic_pmos I_659(.D(I_659_D), .G(I_659_G), .S(I_691_D));
  generic_nmos I_66(.D(I_67_S), .G(I_65_S), .S(VSS));
  generic_nmos I_660(.D(I_660_D), .G(I_661_G), .S(I_692_D));
  generic_pmos I_661(.D(I_661_D), .G(I_661_G), .S(I_693_D));
  generic_nmos I_662(.D(I_759_D), .G(I_727_D), .S(VSS));
  generic_pmos I_663(.D(I_759_D), .G(I_727_D), .S(VDD));
  generic_nmos I_664(.D(VSS), .G(I_633_D), .S(I_763_D));
  generic_pmos I_665(.D(VDD), .G(I_633_D), .S(I_763_D));
  generic_nmos I_666(.D(I_667_D), .G(I_827_D), .S(I_698_D));
  generic_pmos I_667(.D(I_667_D), .G(I_827_D), .S(I_699_D));
  generic_nmos I_668(.D(I_765_D), .G(I_637_D), .S(I_700_D));
  generic_pmos I_669(.D(VDD), .G(I_637_D), .S(I_765_D));
  generic_pmos I_67(.D(I_67_D), .G(I_65_S), .S(I_67_S));
  generic_nmos I_670(.D(I_670_D), .G(I_671_G), .S(VSS));
  generic_pmos I_671(.D(I_671_D), .G(I_671_G), .S(VDD));
  generic_nmos I_672(.D(VSS), .G(I_768_D), .S(I_705_D));
  generic_pmos I_673(.D(VDD), .G(I_768_D), .S(I_705_D));
  generic_nmos I_674(.D(I_674_D), .G(I_1249_D), .S(VSS));
  generic_pmos I_675(.D(I_675_D), .G(I_1249_D), .S(VDD));
  generic_nmos I_676(.D(I_676_D), .G(I_709_S), .S(VSS));
  generic_pmos I_677(.D(I_741_D), .G(I_709_S), .S(VDD));
  generic_nmos I_678(.D(VSS), .G(I_1187_S), .S(I_710_D));
  generic_pmos I_679(.D(VDD), .G(I_1187_S), .S(I_773_S));
  generic_nmos I_68(.D(VSS), .G(I_133_D), .S(I_69_S));
  generic_nmos I_680(.D(I_680_D), .G(I_681_G), .S(VSS));
  generic_pmos I_681(.D(I_681_D), .G(I_681_G), .S(VDD));
  generic_nmos I_682(.D(I_682_D), .G(I_616_S), .S(I_714_D));
  generic_pmos I_683(.D(VDD), .G(I_616_S), .S(I_715_D));
  generic_nmos I_684(.D(I_684_D), .G(I_685_G), .S(I_716_D));
  generic_pmos I_685(.D(I_685_D), .G(I_685_G), .S(I_717_D));
  generic_nmos I_686(.D(I_686_D), .G(I_687_G), .S(I_718_D));
  generic_pmos I_687(.D(I_687_D), .G(I_687_G), .S(I_719_D));
  generic_nmos I_688(.D(I_688_D), .G(I_689_G), .S(I_720_D));
  generic_pmos I_689(.D(I_689_D), .G(I_689_G), .S(I_721_D));
  generic_pmos I_69(.D(VDD), .G(I_133_D), .S(I_69_S));
  generic_nmos I_690(.D(I_690_D), .G(I_691_G), .S(I_722_D));
  generic_pmos I_691(.D(I_691_D), .G(I_691_G), .S(I_723_D));
  generic_nmos I_692(.D(I_692_D), .G(I_693_G), .S(VSS));
  generic_pmos I_693(.D(I_693_D), .G(I_693_G), .S(VDD));
  generic_nmos I_694(.D(VSS), .G(I_791_D), .S(I_727_D));
  generic_pmos I_695(.D(VDD), .G(I_791_D), .S(I_727_D));
  generic_nmos I_696(.D(I_763_D), .G(I_633_D), .S(VSS));
  generic_pmos I_697(.D(I_763_D), .G(I_633_D), .S(VDD));
  generic_nmos I_698(.D(I_698_D), .G(I_827_D), .S(VSS));
  generic_pmos I_699(.D(I_699_D), .G(I_827_D), .S(VDD));
  generic_pmos I_7(.D(I_103_D), .G(I_133_S), .S(VDD));
  generic_nmos I_70(.D(I_70_D), .G(I_135_D), .S(I_133_S));
  generic_nmos I_700(.D(I_700_D), .G(I_799_S), .S(VSS));
  generic_pmos I_701(.D(I_765_D), .G(I_799_S), .S(VDD));
  generic_nmos I_702(.D(VSS), .G(I_575_S), .S(I_735_D));
  generic_pmos I_703(.D(VDD), .G(I_575_S), .S(I_735_D));
  generic_nmos I_704(.D(I_705_D), .G(I_768_D), .S(VSS));
  generic_pmos I_705(.D(I_705_D), .G(I_768_D), .S(VDD));
  generic_nmos I_706(.D(VSS), .G(I_1249_D), .S(I_707_S));
  generic_pmos I_707(.D(VDD), .G(I_1249_D), .S(I_707_S));
  generic_nmos I_708(.D(VSS), .G(I_773_D), .S(I_709_S));
  generic_pmos I_709(.D(VDD), .G(I_773_D), .S(I_709_S));
  generic_pmos I_71(.D(I_133_S), .G(I_135_D), .S(VDD));
  generic_nmos I_710(.D(I_710_D), .G(I_775_D), .S(I_773_S));
  generic_pmos I_711(.D(I_773_S), .G(I_775_D), .S(VDD));
  generic_nmos I_712(.D(VSS), .G(I_235_D), .S(I_713_S));
  generic_pmos I_713(.D(VDD), .G(I_235_D), .S(I_713_S));
  generic_nmos I_714(.D(I_714_D), .G(I_618_S), .S(VSS));
  generic_pmos I_715(.D(I_715_D), .G(I_618_S), .S(VDD));
  generic_nmos I_716(.D(I_716_D), .G(I_717_G), .S(I_716_S));
  generic_pmos I_717(.D(I_717_D), .G(I_717_G), .S(I_717_S));
  generic_nmos I_718(.D(I_718_D), .G(I_719_G), .S(I_718_S));
  generic_pmos I_719(.D(I_719_D), .G(I_719_G), .S(I_719_S));
  generic_nmos I_72(.D(I_72_D), .G(I_73_G), .S(I_72_S));
  generic_nmos I_720(.D(I_720_D), .G(I_721_G), .S(I_720_S));
  generic_pmos I_721(.D(I_721_D), .G(I_721_G), .S(I_721_S));
  generic_nmos I_722(.D(I_722_D), .G(I_723_G), .S(I_722_S));
  generic_pmos I_723(.D(I_723_D), .G(I_723_G), .S(I_723_S));
  generic_nmos I_724(.D(VSS), .G(I_1045_D), .S(I_789_D));
  generic_pmos I_725(.D(VDD), .G(I_1045_D), .S(I_789_D));
  generic_nmos I_726(.D(I_727_D), .G(I_791_D), .S(VSS));
  generic_pmos I_727(.D(I_727_D), .G(I_791_D), .S(VDD));
  generic_nmos I_728(.D(VSS), .G(I_763_D), .S(I_729_S));
  generic_pmos I_729(.D(VDD), .G(I_763_D), .S(I_729_S));
  generic_pmos I_73(.D(I_73_D), .G(I_73_G), .S(I_73_S));
  generic_nmos I_730(.D(VSS), .G(I_731_G), .S(I_730_S));
  generic_pmos I_731(.D(VDD), .G(I_731_G), .S(I_731_S));
  generic_nmos I_732(.D(VSS), .G(I_765_D), .S(I_733_S));
  generic_pmos I_733(.D(VDD), .G(I_765_D), .S(I_733_S));
  generic_nmos I_734(.D(I_735_D), .G(I_575_S), .S(VSS));
  generic_pmos I_735(.D(I_735_D), .G(I_575_S), .S(VDD));
  generic_nmos I_736(.D(VSS), .G(I_865_D), .S(I_768_D));
  generic_pmos I_737(.D(I_768_D), .G(I_1089_D), .S(I_769_D));
  generic_nmos I_738(.D(I_738_D), .G(I_738_G), .S(I_770_D));
  generic_pmos I_739(.D(I_739_D), .G(I_770_G), .S(I_771_D));
  generic_nmos I_74(.D(I_74_D), .G(I_75_G), .S(I_74_S));
  generic_nmos I_740(.D(I_741_D), .G(I_393_S), .S(I_773_D));
  generic_pmos I_741(.D(I_741_D), .G(I_555_D), .S(I_773_D));
  generic_nmos I_742(.D(I_743_D), .G(I_555_D), .S(I_775_D));
  generic_pmos I_743(.D(I_743_D), .G(I_393_S), .S(I_775_D));
  generic_nmos I_744(.D(I_1415_S), .G(I_713_S), .S(I_777_D));
  generic_pmos I_745(.D(I_1415_S), .G(I_779_S), .S(I_777_D));
  generic_nmos I_746(.D(I_779_S), .G(I_713_S), .S(VSS));
  generic_pmos I_747(.D(I_747_D), .G(I_778_G), .S(VDD));
  generic_nmos I_748(.D(I_748_D), .G(I_748_G), .S(I_780_D));
  generic_pmos I_749(.D(I_749_D), .G(I_780_G), .S(I_781_D));
  generic_pmos I_75(.D(I_75_D), .G(I_75_G), .S(I_75_S));
  generic_nmos I_750(.D(I_750_D), .G(I_750_G), .S(I_782_D));
  generic_pmos I_751(.D(I_751_D), .G(I_782_G), .S(I_783_D));
  generic_nmos I_752(.D(I_752_D), .G(I_752_G), .S(I_784_D));
  generic_pmos I_753(.D(I_753_D), .G(I_784_G), .S(I_785_D));
  generic_nmos I_754(.D(I_754_D), .G(I_754_G), .S(I_786_D));
  generic_pmos I_755(.D(I_755_D), .G(I_786_G), .S(I_787_D));
  generic_nmos I_756(.D(VSS), .G(I_1045_D), .S(I_789_D));
  generic_pmos I_757(.D(VDD), .G(I_1045_D), .S(I_789_D));
  generic_nmos I_758(.D(I_759_D), .G(I_315_D), .S(I_791_D));
  generic_pmos I_759(.D(I_759_D), .G(I_251_S), .S(I_791_D));
  generic_nmos I_76(.D(I_76_D), .G(I_77_G), .S(I_76_S));
  generic_nmos I_760(.D(I_795_D), .G(I_315_D), .S(I_793_D));
  generic_pmos I_761(.D(I_795_D), .G(I_251_S), .S(I_793_D));
  generic_nmos I_762(.D(I_763_D), .G(I_789_D), .S(I_795_D));
  generic_pmos I_763(.D(I_763_D), .G(I_1045_D), .S(I_795_D));
  generic_nmos I_764(.D(I_765_D), .G(I_95_D), .S(I_797_D));
  generic_pmos I_765(.D(I_765_D), .G(I_93_S), .S(I_797_D));
  generic_nmos I_766(.D(I_1407_D), .G(I_93_S), .S(I_799_S));
  generic_pmos I_767(.D(I_767_D), .G(I_798_G), .S(I_1407_D));
  generic_nmos I_768(.D(I_768_D), .G(I_1089_D), .S(VSS));
  generic_pmos I_769(.D(I_769_D), .G(I_865_D), .S(VDD));
  generic_pmos I_77(.D(I_77_D), .G(I_77_G), .S(I_77_S));
  generic_nmos I_770(.D(I_770_D), .G(I_770_G), .S(I_770_S));
  generic_pmos I_771(.D(I_771_D), .G(I_771_G), .S(I_771_S));
  generic_nmos I_772(.D(I_773_D), .G(I_555_D), .S(I_773_S));
  generic_pmos I_773(.D(I_773_D), .G(I_393_S), .S(I_773_S));
  generic_nmos I_774(.D(I_775_D), .G(I_393_S), .S(I_2329_D));
  generic_pmos I_775(.D(I_775_D), .G(I_555_D), .S(I_2329_D));
  generic_nmos I_776(.D(I_777_D), .G(I_779_S), .S(I_873_D));
  generic_pmos I_777(.D(I_777_D), .G(I_713_S), .S(I_873_D));
  generic_nmos I_778(.D(VSS), .G(I_778_G), .S(I_778_S));
  generic_pmos I_779(.D(VDD), .G(I_713_S), .S(I_779_S));
  generic_nmos I_78(.D(I_78_D), .G(I_79_G), .S(I_78_S));
  generic_nmos I_780(.D(I_780_D), .G(I_780_G), .S(I_780_S));
  generic_pmos I_781(.D(I_781_D), .G(I_781_G), .S(I_781_S));
  generic_nmos I_782(.D(I_782_D), .G(I_782_G), .S(I_782_S));
  generic_pmos I_783(.D(I_783_D), .G(I_783_G), .S(I_783_S));
  generic_nmos I_784(.D(I_784_D), .G(I_784_G), .S(I_784_S));
  generic_pmos I_785(.D(I_785_D), .G(I_785_G), .S(I_785_S));
  generic_nmos I_786(.D(I_786_D), .G(I_786_G), .S(I_786_S));
  generic_pmos I_787(.D(I_787_D), .G(I_787_G), .S(I_787_S));
  generic_nmos I_788(.D(I_789_D), .G(I_1045_D), .S(VSS));
  generic_pmos I_789(.D(I_789_D), .G(I_1045_D), .S(VDD));
  generic_pmos I_79(.D(I_79_D), .G(I_79_G), .S(I_79_S));
  generic_nmos I_790(.D(I_791_D), .G(I_251_S), .S(I_855_D));
  generic_pmos I_791(.D(I_791_D), .G(I_315_D), .S(I_855_D));
  generic_nmos I_792(.D(I_793_D), .G(I_251_S), .S(I_825_D));
  generic_pmos I_793(.D(I_793_D), .G(I_315_D), .S(I_825_D));
  generic_nmos I_794(.D(I_795_D), .G(I_1045_D), .S(I_2361_D));
  generic_pmos I_795(.D(I_795_D), .G(I_789_D), .S(I_2361_D));
  generic_nmos I_796(.D(I_797_D), .G(I_93_S), .S(I_925_D));
  generic_pmos I_797(.D(I_797_D), .G(I_95_D), .S(I_925_D));
  generic_nmos I_798(.D(I_799_S), .G(I_798_G), .S(I_798_S));
  generic_pmos I_799(.D(I_1407_D), .G(I_95_D), .S(I_799_S));
  generic_nmos I_8(.D(I_8_D), .G(I_9_G), .S(I_40_D));
  generic_nmos I_80(.D(I_80_D), .G(I_81_G), .S(I_80_S));
  generic_nmos I_800(.D(I_864_D), .G(I_1832_D), .S(I_865_D));
  generic_pmos I_801(.D(VDD), .G(I_1832_D), .S(I_833_D));
  generic_nmos I_802(.D(I_802_D), .G(I_803_G), .S(VSS));
  generic_pmos I_803(.D(I_803_D), .G(I_803_G), .S(VDD));
  generic_nmos I_804(.D(I_901_D), .G(I_1187_S), .S(I_836_D));
  generic_pmos I_805(.D(VDD), .G(I_1187_S), .S(I_901_D));
  generic_nmos I_806(.D(I_903_D), .G(I_933_S), .S(VSS));
  generic_pmos I_807(.D(I_903_D), .G(I_933_S), .S(VDD));
  generic_nmos I_808(.D(I_809_D), .G(I_777_D), .S(VSS));
  generic_pmos I_809(.D(I_809_D), .G(I_777_D), .S(VDD));
  generic_pmos I_81(.D(I_81_D), .G(I_81_G), .S(I_81_S));
  generic_nmos I_810(.D(I_810_D), .G(I_811_G), .S(I_842_D));
  generic_pmos I_811(.D(I_811_D), .G(I_811_G), .S(I_843_D));
  generic_nmos I_812(.D(I_812_D), .G(I_813_G), .S(I_844_D));
  generic_pmos I_813(.D(I_813_D), .G(I_813_G), .S(I_845_D));
  generic_nmos I_814(.D(I_814_D), .G(I_815_G), .S(I_846_D));
  generic_pmos I_815(.D(I_815_D), .G(I_815_G), .S(I_847_D));
  generic_nmos I_816(.D(I_816_D), .G(I_817_G), .S(I_848_D));
  generic_pmos I_817(.D(I_817_D), .G(I_817_G), .S(I_849_D));
  generic_nmos I_818(.D(I_818_D), .G(I_819_G), .S(I_850_D));
  generic_pmos I_819(.D(I_819_D), .G(I_819_G), .S(I_851_D));
  generic_nmos I_82(.D(I_82_D), .G(I_83_G), .S(I_82_S));
  generic_nmos I_820(.D(I_821_D), .G(I_917_D), .S(I_852_D));
  generic_pmos I_821(.D(I_821_D), .G(I_917_D), .S(I_853_D));
  generic_nmos I_822(.D(VSS), .G(I_951_D), .S(I_855_D));
  generic_pmos I_823(.D(VDD), .G(I_951_D), .S(I_855_D));
  generic_nmos I_824(.D(I_825_D), .G(I_921_D), .S(VSS));
  generic_pmos I_825(.D(I_825_D), .G(I_921_D), .S(VDD));
  generic_nmos I_826(.D(I_827_D), .G(I_923_D), .S(I_858_D));
  generic_pmos I_827(.D(I_827_D), .G(I_923_D), .S(I_859_D));
  generic_nmos I_828(.D(I_957_S), .G(I_797_D), .S(VSS));
  generic_pmos I_829(.D(I_957_S), .G(I_797_D), .S(VDD));
  generic_pmos I_83(.D(I_83_D), .G(I_83_G), .S(I_83_S));
  generic_nmos I_830(.D(I_1439_S), .G(I_415_S), .S(I_862_D));
  generic_pmos I_831(.D(I_1439_S), .G(I_415_S), .S(VDD));
  generic_nmos I_832(.D(I_865_D), .G(I_867_D), .S(I_864_D));
  generic_pmos I_833(.D(I_833_D), .G(I_867_D), .S(I_865_D));
  generic_nmos I_834(.D(VSS), .G(I_931_D), .S(I_866_D));
  generic_pmos I_835(.D(VDD), .G(I_931_D), .S(I_867_D));
  generic_nmos I_836(.D(I_836_D), .G(I_869_S), .S(VSS));
  generic_pmos I_837(.D(I_901_D), .G(I_869_S), .S(VDD));
  generic_nmos I_838(.D(VSS), .G(I_1187_S), .S(I_870_D));
  generic_pmos I_839(.D(VDD), .G(I_1187_S), .S(I_933_S));
  generic_nmos I_84(.D(VSS), .G(I_85_G), .S(I_2681_D));
  generic_nmos I_840(.D(VSS), .G(I_809_D), .S(I_873_D));
  generic_pmos I_841(.D(VDD), .G(I_809_D), .S(I_873_D));
  generic_nmos I_842(.D(I_842_D), .G(I_843_G), .S(I_874_D));
  generic_pmos I_843(.D(I_843_D), .G(I_843_G), .S(I_875_D));
  generic_nmos I_844(.D(I_844_D), .G(I_845_G), .S(I_876_D));
  generic_pmos I_845(.D(I_845_D), .G(I_845_G), .S(I_877_D));
  generic_nmos I_846(.D(I_846_D), .G(I_847_G), .S(I_878_D));
  generic_pmos I_847(.D(I_847_D), .G(I_847_G), .S(I_879_D));
  generic_nmos I_848(.D(I_848_D), .G(I_849_G), .S(I_880_D));
  generic_pmos I_849(.D(I_849_D), .G(I_849_G), .S(I_881_D));
  generic_pmos I_85(.D(VDD), .G(I_85_G), .S(I_2681_D));
  generic_nmos I_850(.D(I_850_D), .G(I_851_G), .S(I_882_D));
  generic_pmos I_851(.D(I_851_D), .G(I_851_G), .S(I_883_D));
  generic_nmos I_852(.D(I_852_D), .G(I_917_D), .S(VSS));
  generic_pmos I_853(.D(I_853_D), .G(I_917_D), .S(VDD));
  generic_nmos I_854(.D(I_855_D), .G(I_951_D), .S(VSS));
  generic_pmos I_855(.D(I_855_D), .G(I_951_D), .S(VDD));
  generic_nmos I_856(.D(VSS), .G(I_793_D), .S(I_921_D));
  generic_pmos I_857(.D(VDD), .G(I_793_D), .S(I_921_D));
  generic_nmos I_858(.D(I_858_D), .G(I_923_D), .S(VSS));
  generic_pmos I_859(.D(I_859_D), .G(I_923_D), .S(VDD));
  generic_nmos I_86(.D(VSS), .G(I_87_G), .S(I_2361_D));
  generic_nmos I_860(.D(VSS), .G(I_861_G), .S(VSS));
  generic_pmos I_861(.D(VDD), .G(I_861_G), .S(VDD));
  generic_nmos I_862(.D(I_862_D), .G(I_733_S), .S(I_894_D));
  generic_pmos I_863(.D(VDD), .G(I_733_S), .S(I_1439_S));
  generic_nmos I_864(.D(I_864_D), .G(I_929_D), .S(VSS));
  generic_pmos I_865(.D(I_865_D), .G(I_929_D), .S(VDD));
  generic_nmos I_866(.D(I_866_D), .G(I_995_D), .S(I_867_D));
  generic_pmos I_867(.D(I_867_D), .G(I_995_D), .S(VDD));
  generic_nmos I_868(.D(VSS), .G(I_933_D), .S(I_869_S));
  generic_pmos I_869(.D(VDD), .G(I_933_D), .S(I_869_S));
  generic_pmos I_87(.D(VDD), .G(I_87_G), .S(I_2361_D));
  generic_nmos I_870(.D(I_870_D), .G(I_935_D), .S(I_933_S));
  generic_pmos I_871(.D(I_933_S), .G(I_935_D), .S(VDD));
  generic_nmos I_872(.D(I_873_D), .G(I_809_D), .S(VSS));
  generic_pmos I_873(.D(I_873_D), .G(I_809_D), .S(VDD));
  generic_nmos I_874(.D(I_874_D), .G(I_875_G), .S(I_874_S));
  generic_pmos I_875(.D(I_875_D), .G(I_875_G), .S(I_875_S));
  generic_nmos I_876(.D(I_876_D), .G(I_877_G), .S(I_876_S));
  generic_pmos I_877(.D(I_877_D), .G(I_877_G), .S(I_877_S));
  generic_nmos I_878(.D(I_878_D), .G(I_879_G), .S(I_878_S));
  generic_pmos I_879(.D(I_879_D), .G(I_879_G), .S(I_879_S));
  generic_nmos I_88(.D(I_88_D), .G(I_89_G), .S(I_88_S));
  generic_nmos I_880(.D(I_880_D), .G(I_881_G), .S(I_880_S));
  generic_pmos I_881(.D(I_881_D), .G(I_881_G), .S(I_881_S));
  generic_nmos I_882(.D(I_882_D), .G(I_883_G), .S(I_882_S));
  generic_pmos I_883(.D(I_883_D), .G(I_883_G), .S(I_883_S));
  generic_nmos I_884(.D(VSS), .G(I_885_G), .S(I_884_S));
  generic_pmos I_885(.D(VDD), .G(I_885_G), .S(I_885_S));
  generic_nmos I_886(.D(VSS), .G(I_855_D), .S(I_919_D));
  generic_pmos I_887(.D(VDD), .G(I_855_D), .S(I_919_D));
  generic_nmos I_888(.D(I_921_D), .G(I_793_D), .S(VSS));
  generic_pmos I_889(.D(I_921_D), .G(I_793_D), .S(VDD));
  generic_pmos I_89(.D(I_89_D), .G(I_89_G), .S(I_89_S));
  generic_nmos I_890(.D(VSS), .G(I_891_G), .S(I_890_S));
  generic_pmos I_891(.D(VDD), .G(I_891_G), .S(I_891_S));
  generic_nmos I_892(.D(VSS), .G(I_957_S), .S(I_925_D));
  generic_pmos I_893(.D(VDD), .G(I_957_S), .S(I_925_D));
  generic_nmos I_894(.D(I_894_D), .G(I_1055_S), .S(VSS));
  generic_pmos I_895(.D(I_1439_S), .G(I_1055_S), .S(VDD));
  generic_nmos I_896(.D(VSS), .G(I_867_D), .S(I_928_D));
  generic_pmos I_897(.D(VDD), .G(I_1832_D), .S(I_929_D));
  generic_nmos I_898(.D(I_931_D), .G(I_1027_S), .S(I_930_D));
  generic_pmos I_899(.D(VDD), .G(I_869_S), .S(I_931_D));
  generic_pmos I_9(.D(I_9_D), .G(I_9_G), .S(I_41_D));
  generic_nmos I_90(.D(VSS), .G(I_91_G), .S(I_2041_D));
  generic_nmos I_900(.D(I_901_D), .G(I_393_S), .S(I_933_D));
  generic_pmos I_901(.D(I_901_D), .G(I_555_D), .S(I_933_D));
  generic_nmos I_902(.D(I_903_D), .G(I_555_D), .S(I_935_D));
  generic_pmos I_903(.D(I_903_D), .G(I_393_S), .S(I_935_D));
  generic_nmos I_904(.D(I_2329_D), .G(I_713_S), .S(I_937_D));
  generic_pmos I_905(.D(I_2329_D), .G(I_779_S), .S(I_937_D));
  generic_nmos I_906(.D(I_906_D), .G(I_906_G), .S(I_938_D));
  generic_pmos I_907(.D(I_907_D), .G(I_938_G), .S(I_939_D));
  generic_nmos I_908(.D(I_908_D), .G(I_908_G), .S(I_940_D));
  generic_pmos I_909(.D(I_909_D), .G(I_940_G), .S(I_941_D));
  generic_pmos I_91(.D(VDD), .G(I_91_G), .S(I_2041_D));
  generic_nmos I_910(.D(I_910_D), .G(I_910_G), .S(I_942_D));
  generic_pmos I_911(.D(I_911_D), .G(I_942_G), .S(I_943_D));
  generic_nmos I_912(.D(I_912_D), .G(I_912_G), .S(I_944_D));
  generic_pmos I_913(.D(I_913_D), .G(I_944_G), .S(I_945_D));
  generic_nmos I_914(.D(I_914_D), .G(I_914_G), .S(I_946_D));
  generic_pmos I_915(.D(I_915_D), .G(I_946_G), .S(I_947_D));
  generic_nmos I_916(.D(I_917_D), .G(I_1331_D), .S(I_948_D));
  generic_pmos I_917(.D(I_917_D), .G(I_1331_D), .S(I_949_D));
  generic_nmos I_918(.D(I_919_D), .G(I_251_S), .S(I_951_D));
  generic_pmos I_919(.D(I_919_D), .G(I_315_D), .S(I_951_D));
  generic_nmos I_92(.D(VSS), .G(I_503_G), .S(I_93_S));
  generic_nmos I_920(.D(I_921_D), .G(I_251_S), .S(I_953_D));
  generic_pmos I_921(.D(I_921_D), .G(I_315_D), .S(I_953_D));
  generic_nmos I_922(.D(I_923_D), .G(I_989_D), .S(I_954_D));
  generic_pmos I_923(.D(I_923_D), .G(I_989_D), .S(I_955_D));
  generic_nmos I_924(.D(I_925_D), .G(I_735_D), .S(I_957_D));
  generic_pmos I_925(.D(I_925_D), .G(I_989_D), .S(I_957_D));
  generic_nmos I_926(.D(I_1279_D), .G(I_93_S), .S(I_959_D));
  generic_pmos I_927(.D(I_1279_D), .G(I_95_D), .S(I_959_D));
  generic_nmos I_928(.D(I_928_D), .G(I_1832_D), .S(I_929_D));
  generic_pmos I_929(.D(I_929_D), .G(I_867_D), .S(VDD));
  generic_pmos I_93(.D(VDD), .G(I_503_G), .S(I_93_S));
  generic_nmos I_930(.D(I_930_D), .G(I_869_S), .S(VSS));
  generic_pmos I_931(.D(I_931_D), .G(I_1027_S), .S(VDD));
  generic_nmos I_932(.D(I_933_D), .G(I_555_D), .S(I_933_S));
  generic_pmos I_933(.D(I_933_D), .G(I_393_S), .S(I_933_S));
  generic_nmos I_934(.D(I_935_D), .G(I_393_S), .S(I_1415_S));
  generic_pmos I_935(.D(I_935_D), .G(I_555_D), .S(I_1415_S));
  generic_nmos I_936(.D(I_937_D), .G(I_779_S), .S(I_1033_D));
  generic_pmos I_937(.D(I_937_D), .G(I_713_S), .S(I_1033_D));
  generic_nmos I_938(.D(I_938_D), .G(I_938_G), .S(I_938_S));
  generic_pmos I_939(.D(I_939_D), .G(I_939_G), .S(I_939_S));
  generic_nmos I_94(.D(I_95_D), .G(I_95_G), .S(VSS));
  generic_nmos I_940(.D(I_940_D), .G(I_940_G), .S(I_940_S));
  generic_pmos I_941(.D(I_941_D), .G(I_941_G), .S(I_941_S));
  generic_nmos I_942(.D(I_942_D), .G(I_942_G), .S(I_942_S));
  generic_pmos I_943(.D(I_943_D), .G(I_943_G), .S(I_943_S));
  generic_nmos I_944(.D(I_944_D), .G(I_944_G), .S(I_944_S));
  generic_pmos I_945(.D(I_945_D), .G(I_945_G), .S(I_945_S));
  generic_nmos I_946(.D(I_946_D), .G(I_946_G), .S(I_946_S));
  generic_pmos I_947(.D(I_947_D), .G(I_947_G), .S(I_947_S));
  generic_nmos I_948(.D(I_948_D), .G(I_1331_D), .S(VSS));
  generic_pmos I_949(.D(I_949_D), .G(I_1331_D), .S(VDD));
  generic_pmos I_95(.D(I_95_D), .G(I_95_G), .S(VDD));
  generic_nmos I_950(.D(I_951_D), .G(I_315_D), .S(I_1111_D));
  generic_pmos I_951(.D(I_951_D), .G(I_251_S), .S(I_1111_D));
  generic_nmos I_952(.D(I_953_D), .G(I_315_D), .S(I_1049_S));
  generic_pmos I_953(.D(I_953_D), .G(I_251_S), .S(I_1049_S));
  generic_nmos I_954(.D(I_954_D), .G(I_989_D), .S(VSS));
  generic_pmos I_955(.D(I_955_D), .G(I_989_D), .S(VDD));
  generic_nmos I_956(.D(I_957_D), .G(I_989_D), .S(I_957_S));
  generic_pmos I_957(.D(I_957_D), .G(I_735_D), .S(I_957_S));
  generic_nmos I_958(.D(I_959_D), .G(I_95_D), .S(I_1055_S));
  generic_pmos I_959(.D(I_959_D), .G(I_93_S), .S(I_1055_S));
  generic_nmos I_96(.D(VSS), .G(I_225_D), .S(I_128_D));
  generic_nmos I_960(.D(I_960_D), .G(I_961_G), .S(VSS));
  generic_pmos I_961(.D(I_961_D), .G(I_961_G), .S(VDD));
  generic_nmos I_962(.D(I_995_D), .G(I_1349_D), .S(I_994_D));
  generic_pmos I_963(.D(VDD), .G(I_1349_D), .S(I_995_D));
  generic_nmos I_964(.D(I_1061_D), .G(I_1029_D), .S(VSS));
  generic_pmos I_965(.D(I_1061_D), .G(I_1029_D), .S(VDD));
  generic_nmos I_966(.D(I_1063_D), .G(I_1187_S), .S(I_998_D));
  generic_pmos I_967(.D(VDD), .G(I_1187_S), .S(I_1063_D));
  generic_nmos I_968(.D(I_969_D), .G(I_937_D), .S(VSS));
  generic_pmos I_969(.D(I_969_D), .G(I_937_D), .S(VDD));
  generic_pmos I_97(.D(I_128_D), .G(I_1089_D), .S(I_129_D));
  generic_nmos I_970(.D(I_970_D), .G(I_971_G), .S(I_1002_D));
  generic_pmos I_971(.D(I_971_D), .G(I_971_G), .S(I_1003_D));
  generic_nmos I_972(.D(I_972_D), .G(I_973_G), .S(I_1004_D));
  generic_pmos I_973(.D(I_973_D), .G(I_973_G), .S(I_1005_D));
  generic_nmos I_974(.D(I_975_D), .G(I_1997_D), .S(VSS));
  generic_pmos I_975(.D(I_975_D), .G(I_1997_D), .S(VDD));
  generic_nmos I_976(.D(I_976_D), .G(I_977_G), .S(I_1008_D));
  generic_pmos I_977(.D(I_977_D), .G(I_977_G), .S(I_1009_D));
  generic_nmos I_978(.D(I_978_D), .G(I_979_G), .S(I_1010_D));
  generic_pmos I_979(.D(I_979_D), .G(I_979_G), .S(I_1011_D));
  generic_nmos I_98(.D(I_131_S), .G(I_67_S), .S(VSS));
  generic_nmos I_980(.D(I_1045_D), .G(I_983_D), .S(VSS));
  generic_pmos I_981(.D(I_1045_D), .G(I_983_D), .S(VDD));
  generic_nmos I_982(.D(I_983_D), .G(I_1113_S), .S(I_1014_D));
  generic_pmos I_983(.D(I_983_D), .G(I_1113_S), .S(I_1015_D));
  generic_nmos I_984(.D(VSS), .G(I_953_D), .S(I_1401_D));
  generic_pmos I_985(.D(VDD), .G(I_953_D), .S(I_1401_D));
  generic_nmos I_986(.D(I_1051_S), .G(I_445_D), .S(VSS));
  generic_pmos I_987(.D(I_1051_S), .G(I_445_D), .S(VDD));
  generic_nmos I_988(.D(I_989_D), .G(I_511_D), .S(VSS));
  generic_pmos I_989(.D(I_989_D), .G(I_511_D), .S(VDD));
  generic_pmos I_99(.D(I_99_D), .G(I_130_G), .S(VDD));
  generic_nmos I_990(.D(I_1087_D), .G(I_959_D), .S(I_1022_D));
  generic_pmos I_991(.D(VDD), .G(I_959_D), .S(I_1087_D));
  generic_nmos I_992(.D(VSS), .G(I_1025_G), .S(I_1025_D));
  generic_pmos I_993(.D(VDD), .G(I_1025_G), .S(I_1025_D));
  generic_nmos I_994(.D(I_994_D), .G(I_1249_D), .S(VSS));
  generic_pmos I_995(.D(I_995_D), .G(I_1249_D), .S(VDD));
  generic_nmos I_996(.D(VSS), .G(I_1187_S), .S(I_1028_D));
  generic_pmos I_997(.D(VDD), .G(I_1187_S), .S(I_1029_D));
  generic_nmos I_998(.D(I_998_D), .G(I_1093_S), .S(VSS));
  generic_pmos I_999(.D(I_1063_D), .G(I_1093_S), .S(VDD));

  //--------------------------------------------------------------------------
  // Output assignments
  //--------------------------------------------------------------------------

  // Inverting pin drivers
  assign RC0   = !I_3519_D;
  assign RC1   = !I_3675_D;
  assign RC2   = !I_3999_D;
  assign RC3   = !I_1919_D;
  assign RC4   = !I_2399_D;
  assign RC5   = !I_2879_D;
  assign RC6   = !I_3359_D;
  assign RC7   = !I_3423_D;
  assign MXSEL = !I_1757_D;
  assign nROM  = !I_3331_D;

  // Noninverting pin drivers
  assign PHI  = I_245_D;
  assign CAS  = I_59_D;
  assign RAS  = I_821_D;
  assign WE   = I_3979_D;
  assign nIO  = I_3651_D;

  // Video outputs
  // For the inverting output driver of the RED pad:
  // * I_131_S goes to the pmos gate and
  // * I_321_D goes to the nmos gate.
  // Here we use the pmos control, since its behaviour looks more appropriate.
  assign RED   = !I_131_S;
  assign GREEN = !I_385_D;
  assign BLUE  = !I_705_D;
  assign SYNC  = I_3_G;

endmodule
