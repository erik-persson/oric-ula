//----------------------------------------------------------------------------
//
//  CMOS transistor netlist for the Oric HCS10017 ULA, processed version
//
//  Generated from an ULA die photograph in 2018 by Mike Connors, Datel
//  https://www.rawscience.co.uk/
//
//  Originally published by Mike Brown
//  https://oric.signal11.org.uk/html/ula-dieshot.htm
//
//  Re-used in oric-ula project by Erik Persson, 2023
//  https://github.com/erik-persson/oric-ula
//
//----------------------------------------------------------------------------

module Top();
supply1  VDD;
supply0  VSS;
wire  auto_net_1;
wire  auto_net_2;
wire  auto_net_3;
wire  auto_net_4;
wire  I_1002_D;
wire  I_1003_D;
wire  I_1003_G;
wire  I_1004_D;
wire  I_1005_D;
wire  I_1005_G;
wire  I_1008_D;
wire  I_1009_D;
wire  I_1009_G;
wire  I_1010_D;
wire  I_1011_D;
wire  I_1011_G;
wire  I_1014_D;
wire  I_1015_D;
wire  I_1019_G;
wire  I_101_D;
wire  I_1022_D;
wire  I_1025_D;
wire  I_1025_G;
wire  I_1027_S;
wire  I_1028_D;
wire  I_1029_D;
wire  I_1033_D;
wire  I_1034_D;
wire  I_1034_S;
wire  I_1035_D;
wire  I_1035_G;
wire  I_1035_S;
wire  I_1036_D;
wire  I_1036_S;
wire  I_1037_D;
wire  I_1037_G;
wire  I_1037_S;
wire  I_1038_D;
wire  I_1039_D;
wire  I_103_D;
wire  I_1040_D;
wire  I_1040_S;
wire  I_1041_D;
wire  I_1041_G;
wire  I_1041_S;
wire  I_1042_D;
wire  I_1042_S;
wire  I_1043_D;
wire  I_1043_G;
wire  I_1043_S;
wire  I_1045_D;
wire  I_1046_S;
wire  I_1047_G;
wire  I_1047_S;
wire  I_1049_S;
wire  I_104_D;
wire  I_104_G;
wire  I_1051_S;
wire  I_1055_S;
wire  I_105_D;
wire  I_1061_D;
wire  I_1063_D;
wire  I_1065_D;
wire  I_1067_D;
wire  I_1069_D;
wire  I_106_D;
wire  I_106_G;
wire  I_1072_D;
wire  I_1072_G;
wire  I_1073_D;
wire  I_1074_D;
wire  I_1074_G;
wire  I_1075_D;
wire  I_1076_D;
wire  I_1076_G;
wire  I_1077_D;
wire  I_107_D;
wire  I_1085_D;
wire  I_1087_D;
wire  I_1088_D;
wire  I_1089_D;
wire  I_108_D;
wire  I_108_G;
wire  I_1090_D;
wire  I_1091_D;
wire  I_1093_D;
wire  I_1093_S;
wire  I_1095_D;
wire  I_1096_G;
wire  I_1096_S;
wire  I_1097_S;
wire  I_1098_G;
wire  I_1098_S;
wire  I_1099_S;
wire  I_109_D;
wire  I_10_D;
wire  I_1100_G;
wire  I_1100_S;
wire  I_1101_S;
wire  I_1102_D;
wire  I_1103_D;
wire  I_1104_D;
wire  I_1104_G;
wire  I_1104_S;
wire  I_1105_D;
wire  I_1105_G;
wire  I_1105_S;
wire  I_1106_D;
wire  I_1106_G;
wire  I_1106_S;
wire  I_1107_D;
wire  I_1107_G;
wire  I_1107_S;
wire  I_1108_D;
wire  I_1108_G;
wire  I_1108_S;
wire  I_1109_D;
wire  I_1109_G;
wire  I_1109_S;
wire  I_110_D;
wire  I_110_G;
wire  I_1111_D;
wire  I_1112_D;
wire  I_1113_D;
wire  I_1113_S;
wire  I_1114_D;
wire  I_1115_D;
wire  I_1116_G;
wire  I_1116_S;
wire  I_1117_D;
wire  I_1119_D;
wire  I_111_D;
wire  I_1120_D;
wire  I_1121_D;
wire  I_1121_G;
wire  I_112_D;
wire  I_112_G;
wire  I_1132_D;
wire  I_1133_D;
wire  I_1133_G;
wire  I_1136_D;
wire  I_1137_D;
wire  I_1137_G;
wire  I_1139_D;
wire  I_113_D;
wire  I_1144_D;
wire  I_1145_D;
wire  I_1145_G;
wire  I_114_D;
wire  I_114_G;
wire  I_1153_G;
wire  I_1158_D;
wire  I_115_D;
wire  I_1164_D;
wire  I_1165_D;
wire  I_1165_G;
wire  I_1166_D;
wire  I_1168_D;
wire  I_1169_D;
wire  I_1169_G;
wire  I_116_D;
wire  I_116_G;
wire  I_1178_D;
wire  I_117_D;
wire  I_1180_D;
wire  I_1183_G;
wire  I_1184_D;
wire  I_1185_D;
wire  I_1185_G;
wire  I_1187_S;
wire  I_1188_D;
wire  I_1189_D;
wire  I_118_D;
wire  I_118_G;
wire  I_1193_G;
wire  I_1195_D;
wire  I_1196_D;
wire  I_1196_S;
wire  I_1197_D;
wire  I_1197_G;
wire  I_1197_S;
wire  I_1198_S;
wire  I_1199_G;
wire  I_1199_S;
wire  I_11_D;
wire  I_11_G;
wire  I_1200_D;
wire  I_1200_S;
wire  I_1201_D;
wire  I_1201_G;
wire  I_1201_S;
wire  I_1205_D;
wire  I_1207_D;
wire  I_1208_D;
wire  I_1209_D;
wire  I_1209_S;
wire  I_1210_D;
wire  I_1211_D;
wire  I_1212_D;
wire  I_1213_D;
wire  I_1221_D;
wire  I_1223_D;
wire  I_1225_D;
wire  I_1227_D;
wire  I_1228_D;
wire  I_1228_G;
wire  I_1230_D;
wire  I_1230_G;
wire  I_1235_D;
wire  I_1237_D;
wire  I_1239_D;
wire  I_1244_D;
wire  I_1244_G;
wire  I_1247_D;
wire  I_1249_D;
wire  I_1250_D;
wire  I_1250_G;
wire  I_1251_D;
wire  I_1253_D;
wire  I_1253_S;
wire  I_1255_D;
wire  I_1257_D;
wire  I_1258_G;
wire  I_1259_D;
wire  I_1259_S;
wire  I_1260_G;
wire  I_1261_G;
wire  I_1261_S;
wire  I_1262_G;
wire  I_1263_G;
wire  I_1263_S;
wire  I_1265_D;
wire  I_1267_D;
wire  I_1267_S;
wire  I_1269_D;
wire  I_1269_S;
wire  I_1271_D;
wire  I_1272_D;
wire  I_1273_D;
wire  I_1273_S;
wire  I_1274_D;
wire  I_1275_D;
wire  I_1279_D;
wire  I_1279_S;
wire  I_127_D;
wire  I_1280_D;
wire  I_1281_D;
wire  I_1281_G;
wire  I_1283_D;
wire  I_128_D;
wire  I_1292_D;
wire  I_1293_D;
wire  I_1293_G;
wire  I_1295_D;
wire  I_1297_D;
wire  I_1298_D;
wire  I_1299_D;
wire  I_1299_G;
wire  I_129_D;
wire  I_12_D;
wire  I_1301_D;
wire  I_1304_D;
wire  I_1305_D;
wire  I_1305_G;
wire  I_1307_D;
wire  I_1309_D;
wire  I_130_G;
wire  I_130_S;
wire  I_1311_G;
wire  I_1313_G;
wire  I_1318_D;
wire  I_131_S;
wire  I_1324_D;
wire  I_1325_D;
wire  I_1325_G;
wire  I_1329_G;
wire  I_1331_D;
wire  I_1335_D;
wire  I_133_D;
wire  I_133_S;
wire  I_1340_D;
wire  I_1341_D;
wire  I_1342_D;
wire  I_1343_D;
wire  I_1344_D;
wire  I_1345_D;
wire  I_1347_D;
wire  I_1348_D;
wire  I_1349_D;
wire  I_1355_D;
wire  I_1356_D;
wire  I_1356_S;
wire  I_1357_D;
wire  I_1357_G;
wire  I_1357_S;
wire  I_1358_D;
wire  I_1359_D;
wire  I_135_D;
wire  I_1361_S;
wire  I_1362_D;
wire  I_1363_D;
wire  I_1364_D;
wire  I_1365_D;
wire  I_1365_S;
wire  I_1368_D;
wire  I_1369_D;
wire  I_1369_S;
wire  I_136_D;
wire  I_136_G;
wire  I_136_S;
wire  I_1371_D;
wire  I_1373_S;
wire  I_1374_S;
wire  I_1375_G;
wire  I_1375_S;
wire  I_1379_D;
wire  I_137_D;
wire  I_137_G;
wire  I_137_S;
wire  I_1381_D;
wire  I_1383_D;
wire  I_1385_D;
wire  I_1387_D;
wire  I_1388_D;
wire  I_1388_G;
wire  I_138_D;
wire  I_138_G;
wire  I_138_S;
wire  I_1393_D;
wire  I_1397_D;
wire  I_1399_D;
wire  I_139_D;
wire  I_139_G;
wire  I_139_S;
wire  I_13_D;
wire  I_13_G;
wire  I_1401_D;
wire  I_1402_D;
wire  I_1402_G;
wire  I_1403_D;
wire  I_1407_D;
wire  I_1408_D;
wire  I_1408_G;
wire  I_1409_D;
wire  I_1409_G;
wire  I_140_D;
wire  I_140_G;
wire  I_140_S;
wire  I_1410_G;
wire  I_1410_S;
wire  I_1411_S;
wire  I_1413_D;
wire  I_1413_S;
wire  I_1415_D;
wire  I_1415_S;
wire  I_1417_D;
wire  I_1417_S;
wire  I_1419_D;
wire  I_1419_S;
wire  I_141_D;
wire  I_141_G;
wire  I_141_S;
wire  I_1420_S;
wire  I_1421_G;
wire  I_1421_S;
wire  I_1422_D;
wire  I_1423_D;
wire  I_1425_S;
wire  I_1427_D;
wire  I_1429_D;
wire  I_142_D;
wire  I_142_G;
wire  I_142_S;
wire  I_1431_D;
wire  I_1433_D;
wire  I_1435_D;
wire  I_1435_G;
wire  I_1435_S;
wire  I_1437_D;
wire  I_1439_D;
wire  I_1439_S;
wire  I_143_D;
wire  I_143_G;
wire  I_143_S;
wire  I_1448_D;
wire  I_1449_D;
wire  I_1449_G;
wire  I_144_D;
wire  I_144_G;
wire  I_144_S;
wire  I_1452_D;
wire  I_1453_D;
wire  I_1453_G;
wire  I_1456_D;
wire  I_1457_D;
wire  I_1457_G;
wire  I_145_D;
wire  I_145_G;
wire  I_145_S;
wire  I_1461_D;
wire  I_1469_D;
wire  I_146_D;
wire  I_146_G;
wire  I_146_S;
wire  I_1478_D;
wire  I_147_D;
wire  I_147_G;
wire  I_147_S;
wire  I_1480_D;
wire  I_1481_D;
wire  I_1481_G;
wire  I_1482_D;
wire  I_1483_D;
wire  I_1484_D;
wire  I_1485_D;
wire  I_1485_G;
wire  I_1486_D;
wire  I_1488_D;
wire  I_1489_D;
wire  I_1489_G;
wire  I_148_D;
wire  I_148_G;
wire  I_148_S;
wire  I_1491_D;
wire  I_1498_D;
wire  I_1499_D;
wire  I_149_D;
wire  I_149_G;
wire  I_149_S;
wire  I_14_D;
wire  I_1502_D;
wire  I_1507_D;
wire  I_1508_D;
wire  I_1511_S;
wire  I_1512_D;
wire  I_1512_S;
wire  I_1513_D;
wire  I_1513_G;
wire  I_1513_S;
wire  I_1515_S;
wire  I_1516_D;
wire  I_1516_S;
wire  I_1517_D;
wire  I_1517_G;
wire  I_1517_S;
wire  I_1518_D;
wire  I_1518_S;
wire  I_1519_G;
wire  I_1519_S;
wire  I_151_D;
wire  I_151_G;
wire  I_1520_D;
wire  I_1520_S;
wire  I_1521_D;
wire  I_1521_G;
wire  I_1521_S;
wire  I_1523_S;
wire  I_1525_D;
wire  I_1529_D;
wire  I_1531_S;
wire  I_1534_D;
wire  I_1535_D;
wire  I_1537_D;
wire  I_1539_D;
wire  I_153_D;
wire  I_1541_D;
wire  I_1544_D;
wire  I_1544_G;
wire  I_1546_D;
wire  I_1546_G;
wire  I_1547_D;
wire  I_1548_D;
wire  I_1548_G;
wire  I_1549_D;
wire  I_1550_D;
wire  I_1550_G;
wire  I_1551_D;
wire  I_1554_D;
wire  I_1554_G;
wire  I_1555_D;
wire  I_1559_D;
wire  I_155_D;
wire  I_1561_D;
wire  I_1569_D;
wire  I_1571_D;
wire  I_1571_S;
wire  I_1573_D;
wire  I_1573_S;
wire  I_1575_D;
wire  I_1575_S;
wire  I_1576_S;
wire  I_1577_G;
wire  I_1577_S;
wire  I_1578_D;
wire  I_1578_G;
wire  I_1578_S;
wire  I_1579_D;
wire  I_1579_G;
wire  I_1579_S;
wire  I_157_D;
wire  I_1580_D;
wire  I_1580_G;
wire  I_1580_S;
wire  I_1581_D;
wire  I_1581_G;
wire  I_1581_S;
wire  I_1582_D;
wire  I_1582_G;
wire  I_1582_S;
wire  I_1583_D;
wire  I_1583_G;
wire  I_1583_S;
wire  I_1584_D;
wire  I_1585_D;
wire  I_1586_D;
wire  I_1586_G;
wire  I_1586_S;
wire  I_1587_D;
wire  I_1587_G;
wire  I_1587_S;
wire  I_1588_S;
wire  I_1589_S;
wire  I_158_G;
wire  I_158_S;
wire  I_1591_D;
wire  I_1593_D;
wire  I_1593_S;
wire  I_1597_D;
wire  I_1598_S;
wire  I_1599_S;
wire  I_159_S;
wire  I_15_D;
wire  I_15_G;
wire  I_1609_D;
wire  I_1610_D;
wire  I_1611_D;
wire  I_1611_G;
wire  I_1612_D;
wire  I_1613_D;
wire  I_1613_G;
wire  I_1614_D;
wire  I_1615_D;
wire  I_1615_G;
wire  I_1618_D;
wire  I_1619_D;
wire  I_1619_G;
wire  I_1620_D;
wire  I_1621_D;
wire  I_1621_G;
wire  I_1623_D;
wire  I_1627_D;
wire  I_162_D;
wire  I_1631_G;
wire  I_1638_D;
wire  I_163_D;
wire  I_163_G;
wire  I_1642_D;
wire  I_1643_D;
wire  I_1643_G;
wire  I_1644_D;
wire  I_1645_D;
wire  I_1645_G;
wire  I_1648_D;
wire  I_1649_D;
wire  I_1650_D;
wire  I_1651_D;
wire  I_1651_G;
wire  I_1660_D;
wire  I_1662_D;
wire  I_1667_D;
wire  I_1668_D;
wire  I_1671_S;
wire  I_1672_D;
wire  I_1673_D;
wire  I_1674_D;
wire  I_1674_S;
wire  I_1675_D;
wire  I_1675_G;
wire  I_1675_S;
wire  I_1676_D;
wire  I_1676_S;
wire  I_1677_D;
wire  I_1677_G;
wire  I_1677_S;
wire  I_1678_D;
wire  I_1679_D;
wire  I_1681_S;
wire  I_1682_D;
wire  I_1682_S;
wire  I_1683_D;
wire  I_1683_G;
wire  I_1683_S;
wire  I_1684_S;
wire  I_1685_D;
wire  I_1685_G;
wire  I_1685_S;
wire  I_1687_S;
wire  I_1689_D;
wire  I_168_D;
wire  I_1692_D;
wire  I_1693_D;
wire  I_1694_D;
wire  I_1695_D;
wire  I_1697_D;
wire  I_1699_D;
wire  I_169_D;
wire  I_169_G;
wire  I_16_D;
wire  I_1701_D;
wire  I_1706_D;
wire  I_1706_G;
wire  I_1707_D;
wire  I_1709_D;
wire  I_1713_D;
wire  I_1715_D;
wire  I_1729_D;
wire  I_1729_S;
wire  I_172_D;
wire  I_1730_G;
wire  I_1731_D;
wire  I_1731_S;
wire  I_1733_D;
wire  I_1733_S;
wire  I_1735_D;
wire  I_1735_S;
wire  I_1736_D;
wire  I_1737_D;
wire  I_1738_D;
wire  I_1738_G;
wire  I_1738_S;
wire  I_1739_D;
wire  I_1739_G;
wire  I_1739_S;
wire  I_173_D;
wire  I_173_G;
wire  I_1740_G;
wire  I_1740_S;
wire  I_1741_S;
wire  I_1742_D;
wire  I_1743_D;
wire  I_1744_G;
wire  I_1744_S;
wire  I_1746_G;
wire  I_1746_S;
wire  I_1748_S;
wire  I_1749_S;
wire  I_174_D;
wire  I_1750_S;
wire  I_1751_S;
wire  I_1752_S;
wire  I_1753_S;
wire  I_1755_D;
wire  I_1757_D;
wire  I_1758_S;
wire  I_1759_S;
wire  I_175_D;
wire  I_175_G;
wire  I_1761_D;
wire  I_1761_G;
wire  I_1763_D;
wire  I_176_D;
wire  I_1770_D;
wire  I_1771_D;
wire  I_1771_G;
wire  I_1772_D;
wire  I_1773_D;
wire  I_1773_G;
wire  I_1778_D;
wire  I_1779_D;
wire  I_1779_G;
wire  I_177_D;
wire  I_177_G;
wire  I_178_D;
wire  I_1798_D;
wire  I_179_D;
wire  I_179_G;
wire  I_17_D;
wire  I_17_G;
wire  I_1800_D;
wire  I_1802_D;
wire  I_1803_D;
wire  I_1803_G;
wire  I_1804_D;
wire  I_1805_D;
wire  I_1805_G;
wire  I_1806_D;
wire  I_1807_D;
wire  I_1808_D;
wire  I_1810_D;
wire  I_1811_D;
wire  I_1811_G;
wire  I_1812_D;
wire  I_1821_D;
wire  I_1822_D;
wire  I_1825_D;
wire  I_1826_D;
wire  I_1828_D;
wire  I_1831_S;
wire  I_1832_D;
wire  I_1832_S;
wire  I_1833_G;
wire  I_1833_S;
wire  I_1834_D;
wire  I_1834_S;
wire  I_1835_D;
wire  I_1835_G;
wire  I_1835_S;
wire  I_1836_D;
wire  I_1836_S;
wire  I_1837_D;
wire  I_1837_G;
wire  I_1837_S;
wire  I_1839_S;
wire  I_1843_S;
wire  I_1844_D;
wire  I_1845_D;
wire  I_1847_D;
wire  I_1853_S;
wire  I_1854_D;
wire  I_1855_D;
wire  I_1858_D;
wire  I_185_D;
wire  I_1861_D;
wire  I_1864_D;
wire  I_1864_G;
wire  I_1865_D;
wire  I_1870_D;
wire  I_1870_G;
wire  I_1871_D;
wire  I_1873_D;
wire  I_1874_D;
wire  I_1874_G;
wire  I_1876_D;
wire  I_1876_G;
wire  I_1879_D;
wire  I_1881_D;
wire  I_1888_D;
wire  I_1888_G;
wire  I_1889_D;
wire  I_1890_D;
wire  I_1891_S;
wire  I_1893_D;
wire  I_1893_S;
wire  I_1895_D;
wire  I_1895_S;
wire  I_1896_D;
wire  I_1896_G;
wire  I_1896_S;
wire  I_1897_D;
wire  I_1897_G;
wire  I_1897_S;
wire  I_1899_D;
wire  I_1899_S;
wire  I_18_D;
wire  I_1900_D;
wire  I_1901_D;
wire  I_1902_D;
wire  I_1902_G;
wire  I_1902_S;
wire  I_1903_D;
wire  I_1903_G;
wire  I_1903_S;
wire  I_1904_G;
wire  I_1904_S;
wire  I_1906_S;
wire  I_1907_G;
wire  I_1907_S;
wire  I_1908_S;
wire  I_1909_G;
wire  I_1909_S;
wire  I_190_D;
wire  I_1911_D;
wire  I_1911_S;
wire  I_1913_D;
wire  I_1913_S;
wire  I_1915_D;
wire  I_1915_S;
wire  I_1916_D;
wire  I_1917_D;
wire  I_1919_D;
wire  I_191_D;
wire  I_191_G;
wire  I_1921_G;
wire  I_1923_D;
wire  I_1928_D;
wire  I_1929_D;
wire  I_1929_G;
wire  I_1934_D;
wire  I_1935_D;
wire  I_1935_G;
wire  I_1936_D;
wire  I_1937_D;
wire  I_1937_G;
wire  I_1938_D;
wire  I_1939_D;
wire  I_1939_G;
wire  I_193_D;
wire  I_1943_D;
wire  I_1946_D;
wire  I_1947_D;
wire  I_1947_G;
wire  I_1949_D;
wire  I_1952_D;
wire  I_1958_D;
wire  I_1960_D;
wire  I_1961_D;
wire  I_1961_G;
wire  I_1962_D;
wire  I_1969_D;
wire  I_196_D;
wire  I_1970_D;
wire  I_1971_D;
wire  I_1971_G;
wire  I_1973_D;
wire  I_1982_D;
wire  I_1985_S;
wire  I_1986_D;
wire  I_1987_D;
wire  I_1988_D;
wire  I_1991_S;
wire  I_1992_D;
wire  I_1992_S;
wire  I_1993_D;
wire  I_1993_G;
wire  I_1993_S;
wire  I_1994_D;
wire  I_1995_S;
wire  I_1997_D;
wire  I_1998_D;
wire  I_1999_D;
wire  I_19_D;
wire  I_19_G;
wire  I_2001_S;
wire  I_2002_D;
wire  I_2002_S;
wire  I_2003_D;
wire  I_2003_G;
wire  I_2003_S;
wire  I_2004_S;
wire  I_2005_G;
wire  I_2005_S;
wire  I_2007_D;
wire  I_2009_D;
wire  I_200_D;
wire  I_2010_D;
wire  I_2011_D;
wire  I_2012_D;
wire  I_2013_D;
wire  I_2014_D;
wire  I_2015_D;
wire  I_201_D;
wire  I_201_G;
wire  I_2021_D;
wire  I_2024_D;
wire  I_2024_G;
wire  I_2025_D;
wire  I_2026_D;
wire  I_2026_G;
wire  I_2028_D;
wire  I_2028_G;
wire  I_2029_D;
wire  I_202_D;
wire  I_2033_D;
wire  I_2034_D;
wire  I_2034_G;
wire  I_2035_D;
wire  I_2041_D;
wire  I_2049_D;
wire  I_204_D;
wire  I_2050_D;
wire  I_2050_G;
wire  I_2051_D;
wire  I_2053_D;
wire  I_2053_S;
wire  I_2055_D;
wire  I_2055_S;
wire  I_2056_D;
wire  I_2056_G;
wire  I_2056_S;
wire  I_2057_D;
wire  I_2057_G;
wire  I_2057_S;
wire  I_2058_S;
wire  I_2059_G;
wire  I_2059_S;
wire  I_205_D;
wire  I_205_G;
wire  I_2060_D;
wire  I_2060_G;
wire  I_2060_S;
wire  I_2061_D;
wire  I_2061_G;
wire  I_2061_S;
wire  I_2062_D;
wire  I_2062_G;
wire  I_2063_D;
wire  I_2065_S;
wire  I_2066_D;
wire  I_2066_G;
wire  I_2066_S;
wire  I_2067_D;
wire  I_2067_G;
wire  I_2067_S;
wire  I_2068_D;
wire  I_2069_D;
wire  I_206_D;
wire  I_2071_D;
wire  I_2071_S;
wire  I_2073_D;
wire  I_2074_D;
wire  I_2075_D;
wire  I_2076_D;
wire  I_2077_D;
wire  I_2078_S;
wire  I_2079_S;
wire  I_207_D;
wire  I_207_G;
wire  I_2083_G;
wire  I_2088_D;
wire  I_2089_D;
wire  I_2089_G;
wire  I_208_D;
wire  I_2092_D;
wire  I_2093_D;
wire  I_2093_G;
wire  I_2096_D;
wire  I_2097_D;
wire  I_2097_G;
wire  I_2098_D;
wire  I_2099_D;
wire  I_2099_G;
wire  I_209_D;
wire  I_209_G;
wire  I_20_D;
wire  I_2103_D;
wire  I_2105_D;
wire  I_210_D;
wire  I_2112_D;
wire  I_2113_D;
wire  I_2113_G;
wire  I_2114_D;
wire  I_2115_D;
wire  I_2118_D;
wire  I_211_D;
wire  I_211_G;
wire  I_2120_D;
wire  I_2121_D;
wire  I_2121_G;
wire  I_2123_D;
wire  I_2124_D;
wire  I_2125_D;
wire  I_2125_G;
wire  I_2126_D;
wire  I_2127_D;
wire  I_2128_D;
wire  I_2129_D;
wire  I_2129_G;
wire  I_2130_D;
wire  I_2131_D;
wire  I_2131_G;
wire  I_2132_D;
wire  I_2133_D;
wire  I_2133_G;
wire  I_2135_G;
wire  I_2138_D;
wire  I_2139_D;
wire  I_2140_D;
wire  I_2142_D;
wire  I_2147_S;
wire  I_2148_D;
wire  I_2151_S;
wire  I_2152_D;
wire  I_2152_S;
wire  I_2153_D;
wire  I_2153_G;
wire  I_2153_S;
wire  I_2154_D;
wire  I_2155_D;
wire  I_2157_S;
wire  I_2159_S;
wire  I_2160_D;
wire  I_2160_S;
wire  I_2161_D;
wire  I_2161_G;
wire  I_2161_S;
wire  I_2162_D;
wire  I_2162_S;
wire  I_2163_D;
wire  I_2163_G;
wire  I_2163_S;
wire  I_2165_S;
wire  I_2167_S;
wire  I_2169_D;
wire  I_2171_S;
wire  I_2172_D;
wire  I_2173_D;
wire  I_2174_D;
wire  I_2175_D;
wire  I_2177_D;
wire  I_2181_D;
wire  I_2184_D;
wire  I_2184_G;
wire  I_2185_D;
wire  I_2187_D;
wire  I_2190_D;
wire  I_2190_G;
wire  I_2191_D;
wire  I_2194_D;
wire  I_2194_G;
wire  I_2195_D;
wire  I_2197_D;
wire  I_2199_D;
wire  I_21_D;
wire  I_21_G;
wire  I_2201_D;
wire  I_2209_D;
wire  I_2209_S;
wire  I_220_D;
wire  I_2210_D;
wire  I_2211_D;
wire  I_2213_D;
wire  I_2213_S;
wire  I_2215_D;
wire  I_2215_S;
wire  I_2216_D;
wire  I_2216_G;
wire  I_2216_S;
wire  I_2217_D;
wire  I_2217_G;
wire  I_2217_S;
wire  I_2218_G;
wire  I_2218_S;
wire  I_2219_S;
wire  I_2222_D;
wire  I_2222_G;
wire  I_2222_S;
wire  I_2223_D;
wire  I_2223_G;
wire  I_2223_S;
wire  I_2224_D;
wire  I_2225_D;
wire  I_2226_D;
wire  I_2226_G;
wire  I_2226_S;
wire  I_2227_D;
wire  I_2227_G;
wire  I_2227_S;
wire  I_2228_G;
wire  I_2228_S;
wire  I_222_D;
wire  I_2231_D;
wire  I_2231_S;
wire  I_2233_D;
wire  I_2234_D;
wire  I_2235_D;
wire  I_2236_D;
wire  I_2237_D;
wire  I_2238_S;
wire  I_2239_S;
wire  I_223_D;
wire  I_223_G;
wire  I_2241_G;
wire  I_2248_D;
wire  I_2249_D;
wire  I_2249_G;
wire  I_224_D;
wire  I_2253_D;
wire  I_2254_D;
wire  I_2255_D;
wire  I_2255_G;
wire  I_2258_D;
wire  I_2259_D;
wire  I_2259_G;
wire  I_225_D;
wire  I_2263_D;
wire  I_2265_D;
wire  I_2267_D;
wire  I_2269_D;
wire  I_226_D;
wire  I_2272_D;
wire  I_2274_D;
wire  I_2275_D;
wire  I_2278_D;
wire  I_227_D;
wire  I_2280_D;
wire  I_2281_D;
wire  I_2281_G;
wire  I_2282_D;
wire  I_2285_G;
wire  I_2288_D;
wire  I_2289_D;
wire  I_2290_D;
wire  I_2291_D;
wire  I_2291_G;
wire  I_2292_D;
wire  I_2295_G;
wire  I_229_S;
wire  I_2302_D;
wire  I_2305_S;
wire  I_2306_S;
wire  I_2307_G;
wire  I_2307_S;
wire  I_2308_D;
wire  I_230_D;
wire  I_2311_S;
wire  I_2312_D;
wire  I_2312_S;
wire  I_2313_D;
wire  I_2313_G;
wire  I_2313_S;
wire  I_2314_S;
wire  I_2315_G;
wire  I_2315_S;
wire  I_2317_S;
wire  I_2318_D;
wire  I_2319_D;
wire  I_2321_S;
wire  I_2322_D;
wire  I_2322_S;
wire  I_2323_D;
wire  I_2323_G;
wire  I_2323_S;
wire  I_2329_D;
wire  I_232_D;
wire  I_232_S;
wire  I_2330_D;
wire  I_2331_D;
wire  I_2332_D;
wire  I_2333_D;
wire  I_2334_D;
wire  I_2335_D;
wire  I_233_D;
wire  I_233_G;
wire  I_233_S;
wire  I_2341_D;
wire  I_2344_D;
wire  I_2344_G;
wire  I_2345_D;
wire  I_2348_D;
wire  I_2348_G;
wire  I_234_D;
wire  I_2353_D;
wire  I_2354_D;
wire  I_2354_G;
wire  I_2355_D;
wire  I_2357_D;
wire  I_235_D;
wire  I_2361_D;
wire  I_2369_D;
wire  I_236_D;
wire  I_236_S;
wire  I_2370_G;
wire  I_2371_D;
wire  I_2371_S;
wire  I_2373_D;
wire  I_2373_S;
wire  I_2375_D;
wire  I_2375_S;
wire  I_2376_D;
wire  I_2376_G;
wire  I_2376_S;
wire  I_2377_D;
wire  I_2377_G;
wire  I_2377_S;
wire  I_2379_D;
wire  I_2379_S;
wire  I_237_D;
wire  I_237_G;
wire  I_237_S;
wire  I_2381_G;
wire  I_2381_S;
wire  I_2382_D;
wire  I_2383_D;
wire  I_2384_G;
wire  I_2384_S;
wire  I_2386_D;
wire  I_2386_G;
wire  I_2386_S;
wire  I_2387_D;
wire  I_2387_G;
wire  I_2387_S;
wire  I_2388_G;
wire  I_2388_S;
wire  I_2389_S;
wire  I_238_D;
wire  I_238_S;
wire  I_2390_D;
wire  I_2391_D;
wire  I_2393_D;
wire  I_2394_D;
wire  I_2395_D;
wire  I_2396_D;
wire  I_2397_D;
wire  I_2399_D;
wire  I_239_D;
wire  I_239_G;
wire  I_239_S;
wire  I_23_G;
wire  I_2402_D;
wire  I_2403_D;
wire  I_2403_G;
wire  I_2408_D;
wire  I_2409_D;
wire  I_2409_G;
wire  I_240_D;
wire  I_240_S;
wire  I_2410_D;
wire  I_2411_D;
wire  I_2411_G;
wire  I_2412_D;
wire  I_2413_D;
wire  I_2413_G;
wire  I_2418_D;
wire  I_2419_D;
wire  I_2419_G;
wire  I_241_D;
wire  I_241_G;
wire  I_241_S;
wire  I_2420_D;
wire  I_2421_D;
wire  I_2421_G;
wire  I_2425_D;
wire  I_2427_D;
wire  I_2429_D;
wire  I_242_D;
wire  I_242_S;
wire  I_2432_D;
wire  I_2433_D;
wire  I_2433_G;
wire  I_2434_D;
wire  I_2435_D;
wire  I_2435_G;
wire  I_2438_D;
wire  I_243_D;
wire  I_243_G;
wire  I_243_S;
wire  I_2440_D;
wire  I_2441_D;
wire  I_2441_G;
wire  I_2442_D;
wire  I_2443_D;
wire  I_2443_G;
wire  I_2444_D;
wire  I_2445_D;
wire  I_2445_G;
wire  I_2446_D;
wire  I_2447_D;
wire  I_2448_D;
wire  I_2450_D;
wire  I_2451_D;
wire  I_2451_G;
wire  I_2453_D;
wire  I_2454_D;
wire  I_2455_D;
wire  I_245_D;
wire  I_2462_D;
wire  I_2466_D;
wire  I_2466_S;
wire  I_2467_D;
wire  I_2467_G;
wire  I_2467_S;
wire  I_2468_D;
wire  I_2471_S;
wire  I_2472_D;
wire  I_2472_S;
wire  I_2473_D;
wire  I_2473_G;
wire  I_2473_S;
wire  I_2474_D;
wire  I_2474_S;
wire  I_2475_D;
wire  I_2475_G;
wire  I_2475_S;
wire  I_2476_D;
wire  I_2476_S;
wire  I_2477_D;
wire  I_2477_G;
wire  I_2477_S;
wire  I_2479_S;
wire  I_247_D;
wire  I_2482_D;
wire  I_2482_S;
wire  I_2483_D;
wire  I_2483_G;
wire  I_2483_S;
wire  I_2485_S;
wire  I_2487_S;
wire  I_2489_D;
wire  I_2490_D;
wire  I_2491_D;
wire  I_2492_D;
wire  I_2493_D;
wire  I_2494_D;
wire  I_2495_D;
wire  I_2497_D;
wire  I_2498_D;
wire  I_2498_G;
wire  I_24_D;
wire  I_2501_D;
wire  I_2504_D;
wire  I_2504_G;
wire  I_2505_D;
wire  I_2509_D;
wire  I_2510_D;
wire  I_2510_G;
wire  I_2511_D;
wire  I_2513_D;
wire  I_2514_D;
wire  I_2514_G;
wire  I_2515_D;
wire  I_2517_D;
wire  I_2519_D;
wire  I_251_S;
wire  I_2521_D;
wire  I_2529_D;
wire  I_2529_S;
wire  I_2530_S;
wire  I_2531_G;
wire  I_2531_S;
wire  I_2533_D;
wire  I_2533_S;
wire  I_2534_G;
wire  I_2535_D;
wire  I_2535_G;
wire  I_2535_S;
wire  I_2536_D;
wire  I_2536_G;
wire  I_2536_S;
wire  I_2537_D;
wire  I_2537_G;
wire  I_2537_S;
wire  I_2539_D;
wire  I_2539_S;
wire  I_253_S;
wire  I_2540_G;
wire  I_2540_S;
wire  I_2542_D;
wire  I_2542_G;
wire  I_2542_S;
wire  I_2543_D;
wire  I_2543_G;
wire  I_2543_S;
wire  I_2544_G;
wire  I_2544_S;
wire  I_2545_S;
wire  I_2546_D;
wire  I_2546_G;
wire  I_2546_S;
wire  I_2547_D;
wire  I_2547_G;
wire  I_2547_S;
wire  I_2549_D;
wire  I_2549_S;
wire  I_254_D;
wire  I_254_S;
wire  I_2550_G;
wire  I_2550_S;
wire  I_2553_D;
wire  I_2554_D;
wire  I_2555_D;
wire  I_2556_D;
wire  I_2557_D;
wire  I_2558_S;
wire  I_2559_S;
wire  I_255_D;
wire  I_255_G;
wire  I_255_S;
wire  I_2561_G;
wire  I_2562_D;
wire  I_2563_D;
wire  I_2563_G;
wire  I_2572_D;
wire  I_2573_D;
wire  I_2573_G;
wire  I_2574_D;
wire  I_2575_D;
wire  I_2575_G;
wire  I_2576_D;
wire  I_2577_D;
wire  I_2577_G;
wire  I_2578_D;
wire  I_2579_D;
wire  I_2579_G;
wire  I_2580_D;
wire  I_2581_D;
wire  I_2581_G;
wire  I_2585_D;
wire  I_2592_D;
wire  I_2594_D;
wire  I_2595_D;
wire  I_2595_G;
wire  I_2598_D;
wire  I_25_D;
wire  I_25_G;
wire  I_2601_D;
wire  I_2603_D;
wire  I_2604_D;
wire  I_2605_D;
wire  I_2605_G;
wire  I_2606_D;
wire  I_2607_D;
wire  I_2607_G;
wire  I_2609_D;
wire  I_2610_D;
wire  I_2611_D;
wire  I_2611_G;
wire  I_2612_D;
wire  I_2613_D;
wire  I_2613_G;
wire  I_2614_D;
wire  I_2618_D;
wire  I_261_D;
wire  I_2620_D;
wire  I_2622_D;
wire  I_2625_S;
wire  I_2626_D;
wire  I_2626_S;
wire  I_2627_D;
wire  I_2627_G;
wire  I_2627_S;
wire  I_2628_D;
wire  I_2631_S;
wire  I_2632_D;
wire  I_2633_D;
wire  I_2634_D;
wire  I_2635_D;
wire  I_2636_D;
wire  I_2636_S;
wire  I_2637_D;
wire  I_2637_G;
wire  I_2637_S;
wire  I_2638_D;
wire  I_2638_S;
wire  I_2639_D;
wire  I_2639_G;
wire  I_2639_S;
wire  I_263_D;
wire  I_2641_S;
wire  I_2642_D;
wire  I_2642_S;
wire  I_2643_D;
wire  I_2643_G;
wire  I_2643_S;
wire  I_2644_D;
wire  I_2644_S;
wire  I_2645_D;
wire  I_2645_G;
wire  I_2645_S;
wire  I_2649_D;
wire  I_2650_D;
wire  I_2650_S;
wire  I_2651_G;
wire  I_2651_S;
wire  I_2652_D;
wire  I_2653_D;
wire  I_2654_D;
wire  I_2655_D;
wire  I_2657_D;
wire  I_2658_D;
wire  I_2658_G;
wire  I_2659_D;
wire  I_265_D;
wire  I_2661_D;
wire  I_2664_D;
wire  I_2664_G;
wire  I_2665_D;
wire  I_2668_D;
wire  I_2668_G;
wire  I_2669_D;
wire  I_266_D;
wire  I_266_G;
wire  I_2673_D;
wire  I_2674_D;
wire  I_2674_G;
wire  I_2675_D;
wire  I_2679_D;
wire  I_267_D;
wire  I_2681_D;
wire  I_2689_D;
wire  I_268_D;
wire  I_268_G;
wire  I_2690_D;
wire  I_2690_G;
wire  I_2690_S;
wire  I_2691_D;
wire  I_2691_G;
wire  I_2691_S;
wire  I_2693_D;
wire  I_2693_S;
wire  I_2695_D;
wire  I_2695_S;
wire  I_2696_D;
wire  I_2696_G;
wire  I_2696_S;
wire  I_2697_D;
wire  I_2697_G;
wire  I_2697_S;
wire  I_2698_D;
wire  I_2699_D;
wire  I_269_D;
wire  I_2700_D;
wire  I_2700_G;
wire  I_2700_S;
wire  I_2701_D;
wire  I_2701_G;
wire  I_2701_S;
wire  I_2705_S;
wire  I_2706_D;
wire  I_2706_G;
wire  I_2706_S;
wire  I_2707_D;
wire  I_2707_G;
wire  I_2707_S;
wire  I_2709_D;
wire  I_2709_S;
wire  I_270_D;
wire  I_270_G;
wire  I_2710_G;
wire  I_2710_S;
wire  I_2711_S;
wire  I_2713_D;
wire  I_2714_D;
wire  I_2715_D;
wire  I_2716_D;
wire  I_2717_D;
wire  I_2718_S;
wire  I_2719_S;
wire  I_271_D;
wire  I_2722_D;
wire  I_2723_D;
wire  I_2723_G;
wire  I_2728_D;
wire  I_2729_D;
wire  I_2729_G;
wire  I_272_D;
wire  I_272_G;
wire  I_2732_D;
wire  I_2733_D;
wire  I_2733_G;
wire  I_2735_D;
wire  I_2736_D;
wire  I_2737_D;
wire  I_2737_G;
wire  I_2738_D;
wire  I_2739_D;
wire  I_2739_G;
wire  I_273_D;
wire  I_2741_D;
wire  I_2742_D;
wire  I_2743_D;
wire  I_2743_G;
wire  I_2745_D;
wire  I_2747_D;
wire  I_2749_D;
wire  I_274_D;
wire  I_274_G;
wire  I_2752_D;
wire  I_2753_D;
wire  I_2753_G;
wire  I_2754_D;
wire  I_2755_D;
wire  I_2755_G;
wire  I_2758_D;
wire  I_275_D;
wire  I_2760_D;
wire  I_2761_D;
wire  I_2761_G;
wire  I_2763_D;
wire  I_2764_D;
wire  I_2765_D;
wire  I_2765_G;
wire  I_2767_G;
wire  I_2770_D;
wire  I_2771_D;
wire  I_2771_G;
wire  I_2773_G;
wire  I_2775_D;
wire  I_277_D;
wire  I_2782_D;
wire  I_2786_D;
wire  I_2786_S;
wire  I_2787_D;
wire  I_2787_G;
wire  I_2787_S;
wire  I_2788_D;
wire  I_2791_S;
wire  I_2792_D;
wire  I_2792_S;
wire  I_2793_D;
wire  I_2793_G;
wire  I_2793_S;
wire  I_2794_D;
wire  I_2795_D;
wire  I_2796_D;
wire  I_2796_S;
wire  I_2797_D;
wire  I_2797_G;
wire  I_2797_S;
wire  I_2799_S;
wire  I_279_D;
wire  I_2800_S;
wire  I_2801_G;
wire  I_2801_S;
wire  I_2805_S;
wire  I_2807_S;
wire  I_2809_D;
wire  I_2810_D;
wire  I_2811_D;
wire  I_2812_D;
wire  I_2813_D;
wire  I_2814_D;
wire  I_2815_D;
wire  I_2817_D;
wire  I_2818_D;
wire  I_2818_G;
wire  I_2819_D;
wire  I_281_D;
wire  I_2821_D;
wire  I_2824_D;
wire  I_2824_G;
wire  I_2825_D;
wire  I_2826_D;
wire  I_2826_G;
wire  I_2828_D;
wire  I_2828_G;
wire  I_2829_D;
wire  I_2830_D;
wire  I_2830_G;
wire  I_2831_D;
wire  I_2834_D;
wire  I_2834_G;
wire  I_2835_D;
wire  I_2837_D;
wire  I_2839_D;
wire  I_2841_D;
wire  I_2849_D;
wire  I_2849_S;
wire  I_2850_D;
wire  I_2850_G;
wire  I_2850_S;
wire  I_2851_D;
wire  I_2851_G;
wire  I_2851_S;
wire  I_2853_D;
wire  I_2853_S;
wire  I_2855_D;
wire  I_2855_S;
wire  I_2856_D;
wire  I_2856_G;
wire  I_2856_S;
wire  I_2857_D;
wire  I_2857_G;
wire  I_2857_S;
wire  I_2859_G;
wire  I_2859_S;
wire  I_285_D;
wire  I_2860_D;
wire  I_2860_G;
wire  I_2860_S;
wire  I_2861_D;
wire  I_2861_G;
wire  I_2861_S;
wire  I_2862_D;
wire  I_2862_G;
wire  I_2862_S;
wire  I_2863_D;
wire  I_2863_G;
wire  I_2863_S;
wire  I_2864_D;
wire  I_2865_D;
wire  I_2866_D;
wire  I_2866_G;
wire  I_2866_S;
wire  I_2867_D;
wire  I_2867_G;
wire  I_2867_S;
wire  I_2869_D;
wire  I_2871_D;
wire  I_2871_S;
wire  I_2873_D;
wire  I_2874_D;
wire  I_2875_D;
wire  I_2876_D;
wire  I_2877_D;
wire  I_2879_D;
wire  I_2881_G;
wire  I_2882_D;
wire  I_2883_D;
wire  I_2883_G;
wire  I_2889_D;
wire  I_288_D;
wire  I_2890_D;
wire  I_2893_D;
wire  I_2894_D;
wire  I_2895_D;
wire  I_2895_G;
wire  I_2898_D;
wire  I_2899_D;
wire  I_2899_G;
wire  I_289_D;
wire  I_2900_D;
wire  I_2901_D;
wire  I_2901_G;
wire  I_2902_D;
wire  I_2903_D;
wire  I_2903_G;
wire  I_2905_D;
wire  I_2907_D;
wire  I_290_D;
wire  I_2912_D;
wire  I_2914_D;
wire  I_2915_D;
wire  I_2915_G;
wire  I_2918_D;
wire  I_291_D;
wire  I_2922_D;
wire  I_2928_D;
wire  I_2929_D;
wire  I_2930_D;
wire  I_2931_D;
wire  I_2931_G;
wire  I_2932_D;
wire  I_2933_D;
wire  I_2933_G;
wire  I_2934_D;
wire  I_2935_D;
wire  I_2935_G;
wire  I_293_D;
wire  I_293_S;
wire  I_2940_D;
wire  I_2942_D;
wire  I_2945_S;
wire  I_2946_D;
wire  I_2946_S;
wire  I_2947_D;
wire  I_2947_G;
wire  I_2947_S;
wire  I_2948_D;
wire  I_2951_S;
wire  I_2952_D;
wire  I_2953_D;
wire  I_2954_D;
wire  I_2955_D;
wire  I_2956_D;
wire  I_2957_D;
wire  I_2958_S;
wire  I_2959_G;
wire  I_2959_S;
wire  I_295_D;
wire  I_2961_S;
wire  I_2962_D;
wire  I_2962_S;
wire  I_2963_D;
wire  I_2963_G;
wire  I_2963_S;
wire  I_2964_D;
wire  I_2964_S;
wire  I_2965_D;
wire  I_2965_G;
wire  I_2965_S;
wire  I_2966_D;
wire  I_2966_S;
wire  I_2967_D;
wire  I_2967_G;
wire  I_2967_S;
wire  I_2969_D;
wire  I_296_G;
wire  I_296_S;
wire  I_2970_D;
wire  I_2971_D;
wire  I_2972_D;
wire  I_2972_S;
wire  I_2973_G;
wire  I_2973_S;
wire  I_2974_D;
wire  I_2975_D;
wire  I_297_S;
wire  I_2981_D;
wire  I_2987_D;
wire  I_298_D;
wire  I_298_G;
wire  I_298_S;
wire  I_2993_D;
wire  I_299_D;
wire  I_299_G;
wire  I_299_S;
wire  I_3004_D;
wire  I_3004_G;
wire  I_3009_D;
wire  I_300_D;
wire  I_300_G;
wire  I_300_S;
wire  I_3010_D;
wire  I_3013_D;
wire  I_3013_S;
wire  I_3015_D;
wire  I_3015_S;
wire  I_3016_D;
wire  I_3017_D;
wire  I_3018_G;
wire  I_3018_S;
wire  I_3019_G;
wire  I_3019_S;
wire  I_301_D;
wire  I_301_G;
wire  I_301_S;
wire  I_3020_D;
wire  I_3021_D;
wire  I_3022_D;
wire  I_3023_D;
wire  I_3024_G;
wire  I_3024_S;
wire  I_3027_D;
wire  I_3029_D;
wire  I_302_D;
wire  I_302_G;
wire  I_302_S;
wire  I_3031_D;
wire  I_3031_S;
wire  I_3033_D;
wire  I_3034_D;
wire  I_3035_D;
wire  I_3036_G;
wire  I_3036_S;
wire  I_3037_G;
wire  I_3037_S;
wire  I_3038_S;
wire  I_3039_S;
wire  I_303_D;
wire  I_303_G;
wire  I_303_S;
wire  I_3042_D;
wire  I_304_D;
wire  I_304_G;
wire  I_304_S;
wire  I_3059_D;
wire  I_305_D;
wire  I_305_G;
wire  I_305_S;
wire  I_3061_D;
wire  I_3063_D;
wire  I_3065_D;
wire  I_306_D;
wire  I_306_G;
wire  I_306_S;
wire  I_3072_D;
wire  I_3073_D;
wire  I_3073_G;
wire  I_3074_D;
wire  I_3075_D;
wire  I_3078_D;
wire  I_307_D;
wire  I_307_G;
wire  I_307_S;
wire  I_3080_D;
wire  I_3082_D;
wire  I_3083_D;
wire  I_3084_D;
wire  I_3086_D;
wire  I_3087_D;
wire  I_3088_D;
wire  I_308_D;
wire  I_3091_G;
wire  I_3093_G;
wire  I_3095_G;
wire  I_3098_D;
wire  I_309_D;
wire  I_3100_D;
wire  I_3102_D;
wire  I_3106_S;
wire  I_3107_G;
wire  I_3107_S;
wire  I_3108_D;
wire  I_3111_S;
wire  I_3112_D;
wire  I_3112_S;
wire  I_3113_G;
wire  I_3113_S;
wire  I_3114_S;
wire  I_3115_G;
wire  I_3115_S;
wire  I_3116_D;
wire  I_3116_S;
wire  I_3117_G;
wire  I_3117_S;
wire  I_3119_S;
wire  I_311_D;
wire  I_3123_S;
wire  I_3125_S;
wire  I_3127_S;
wire  I_3129_D;
wire  I_3130_D;
wire  I_3130_S;
wire  I_3131_G;
wire  I_3131_S;
wire  I_3132_D;
wire  I_3133_D;
wire  I_3134_D;
wire  I_3135_D;
wire  I_3137_D;
wire  I_313_D;
wire  I_3141_D;
wire  I_3146_D;
wire  I_3146_G;
wire  I_3147_D;
wire  I_3148_D;
wire  I_3148_G;
wire  I_3149_D;
wire  I_3151_D;
wire  I_3153_D;
wire  I_3155_D;
wire  I_3157_D;
wire  I_3159_D;
wire  I_315_D;
wire  I_3163_D;
wire  I_3169_D;
wire  I_3169_S;
wire  I_3170_D;
wire  I_3171_D;
wire  I_3173_D;
wire  I_3173_S;
wire  I_3175_D;
wire  I_3175_S;
wire  I_3176_D;
wire  I_3177_D;
wire  I_3178_D;
wire  I_3178_G;
wire  I_3178_S;
wire  I_3179_D;
wire  I_3179_G;
wire  I_3179_S;
wire  I_317_D;
wire  I_3180_D;
wire  I_3180_S;
wire  I_3181_D;
wire  I_3181_G;
wire  I_3181_S;
wire  I_3182_G;
wire  I_3182_S;
wire  I_3184_G;
wire  I_3184_S;
wire  I_3185_S;
wire  I_3189_S;
wire  I_3191_D;
wire  I_3191_S;
wire  I_3192_D;
wire  I_3193_D;
wire  I_3194_G;
wire  I_3194_S;
wire  I_3195_G;
wire  I_3195_S;
wire  I_3196_D;
wire  I_3197_D;
wire  I_3198_S;
wire  I_3199_S;
wire  I_319_D;
wire  I_3201_G;
wire  I_3202_D;
wire  I_3203_D;
wire  I_3203_G;
wire  I_3210_D;
wire  I_3211_D;
wire  I_3211_G;
wire  I_3212_D;
wire  I_3213_D;
wire  I_3213_G;
wire  I_3216_D;
wire  I_3217_D;
wire  I_3217_G;
wire  I_3219_D;
wire  I_321_D;
wire  I_3220_D;
wire  I_3221_D;
wire  I_3221_G;
wire  I_3225_D;
wire  I_3229_D;
wire  I_3232_D;
wire  I_3234_D;
wire  I_3235_D;
wire  I_3235_G;
wire  I_3238_D;
wire  I_3241_D;
wire  I_3242_D;
wire  I_3243_D;
wire  I_3243_G;
wire  I_3244_D;
wire  I_3245_D;
wire  I_3245_G;
wire  I_3246_D;
wire  I_3249_D;
wire  I_3251_G;
wire  I_3254_D;
wire  I_3258_D;
wire  I_3262_D;
wire  I_3265_S;
wire  I_3266_D;
wire  I_3266_S;
wire  I_3267_D;
wire  I_3267_G;
wire  I_3267_S;
wire  I_3268_D;
wire  I_3271_S;
wire  I_3276_D;
wire  I_3276_S;
wire  I_3277_D;
wire  I_3277_G;
wire  I_3277_S;
wire  I_3281_S;
wire  I_3283_S;
wire  I_3284_D;
wire  I_3285_D;
wire  I_3286_D;
wire  I_3287_D;
wire  I_3288_D;
wire  I_3289_D;
wire  I_3290_D;
wire  I_3291_D;
wire  I_3292_D;
wire  I_3293_D;
wire  I_3294_D;
wire  I_3295_D;
wire  I_329_D;
wire  I_32_D;
wire  I_3301_D;
wire  I_3308_D;
wire  I_3308_G;
wire  I_3309_D;
wire  I_3311_D;
wire  I_3313_D;
wire  I_3329_D;
wire  I_332_D;
wire  I_3331_D;
wire  I_3331_G;
wire  I_3333_D;
wire  I_3333_S;
wire  I_3335_D;
wire  I_3335_S;
wire  I_3337_D;
wire  I_3339_D;
wire  I_333_D;
wire  I_333_G;
wire  I_3340_D;
wire  I_3340_G;
wire  I_3340_S;
wire  I_3341_D;
wire  I_3341_G;
wire  I_3341_S;
wire  I_3342_G;
wire  I_3342_S;
wire  I_3345_D;
wire  I_3345_S;
wire  I_3347_D;
wire  I_3348_D;
wire  I_3349_D;
wire  I_334_D;
wire  I_3350_S;
wire  I_3351_S;
wire  I_3352_D;
wire  I_3353_D;
wire  I_3354_S;
wire  I_3355_S;
wire  I_3356_D;
wire  I_3357_D;
wire  I_3359_D;
wire  I_335_D;
wire  I_335_G;
wire  I_3363_D;
wire  I_3369_D;
wire  I_336_D;
wire  I_3371_D;
wire  I_3374_D;
wire  I_3375_D;
wire  I_3375_G;
wire  I_3376_D;
wire  I_3377_D;
wire  I_3377_G;
wire  I_3379_D;
wire  I_337_D;
wire  I_337_G;
wire  I_3381_G;
wire  I_338_D;
wire  I_3392_D;
wire  I_3393_D;
wire  I_3393_G;
wire  I_3398_D;
wire  I_339_D;
wire  I_339_G;
wire  I_33_D;
wire  I_3401_G;
wire  I_3403_G;
wire  I_3407_D;
wire  I_3408_D;
wire  I_3409_D;
wire  I_3409_G;
wire  I_3411_G;
wire  I_3412_D;
wire  I_3413_D;
wire  I_3414_D;
wire  I_3416_D;
wire  I_3418_D;
wire  I_341_D;
wire  I_3420_D;
wire  I_3423_D;
wire  I_3426_D;
wire  I_3427_D;
wire  I_3428_D;
wire  I_3431_S;
wire  I_3433_S;
wire  I_3435_S;
wire  I_3436_D;
wire  I_3439_S;
wire  I_3440_D;
wire  I_3440_S;
wire  I_3441_D;
wire  I_3441_G;
wire  I_3441_S;
wire  I_3443_S;
wire  I_3445_S;
wire  I_3446_D;
wire  I_3447_D;
wire  I_3448_D;
wire  I_3449_D;
wire  I_3450_D;
wire  I_3451_D;
wire  I_3452_D;
wire  I_3453_D;
wire  I_3454_S;
wire  I_3455_G;
wire  I_3455_S;
wire  I_3457_D;
wire  I_3461_D;
wire  I_3465_D;
wire  I_3467_D;
wire  I_3471_D;
wire  I_3475_D;
wire  I_3476_D;
wire  I_3476_G;
wire  I_3477_D;
wire  I_347_D;
wire  I_3480_D;
wire  I_3480_G;
wire  I_3481_D;
wire  I_3489_D;
wire  I_3489_S;
wire  I_3491_D;
wire  I_3491_S;
wire  I_3493_D;
wire  I_3493_S;
wire  I_3495_D;
wire  I_3495_S;
wire  I_3497_S;
wire  I_3499_D;
wire  I_3499_S;
wire  I_3500_D;
wire  I_3501_D;
wire  I_3503_D;
wire  I_3503_S;
wire  I_3504_D;
wire  I_3505_D;
wire  I_3507_D;
wire  I_3508_D;
wire  I_3508_G;
wire  I_3508_S;
wire  I_3509_D;
wire  I_3509_G;
wire  I_3509_S;
wire  I_3510_S;
wire  I_3511_S;
wire  I_3512_D;
wire  I_3512_G;
wire  I_3512_S;
wire  I_3513_D;
wire  I_3513_G;
wire  I_3513_S;
wire  I_3514_S;
wire  I_3515_S;
wire  I_3516_D;
wire  I_3517_D;
wire  I_3519_D;
wire  I_3521_D;
wire  I_3529_D;
wire  I_3529_G;
wire  I_3535_D;
wire  I_3538_D;
wire  I_3539_D;
wire  I_3539_G;
wire  I_3540_D;
wire  I_3541_D;
wire  I_3541_G;
wire  I_3549_D;
wire  I_354_D;
wire  I_3554_D;
wire  I_3555_G;
wire  I_3558_D;
wire  I_355_D;
wire  I_3561_G;
wire  I_3562_D;
wire  I_3563_D;
wire  I_3564_D;
wire  I_3565_D;
wire  I_3567_G;
wire  I_3568_D;
wire  I_3569_D;
wire  I_356_D;
wire  I_3570_D;
wire  I_3571_D;
wire  I_3571_G;
wire  I_3572_D;
wire  I_3573_D;
wire  I_3573_G;
wire  I_3574_D;
wire  I_3576_D;
wire  I_3578_D;
wire  I_3582_D;
wire  I_3584_D;
wire  I_3585_D;
wire  I_3586_D;
wire  I_3587_D;
wire  I_3588_D;
wire  I_3591_S;
wire  I_3593_G;
wire  I_3593_S;
wire  I_3595_S;
wire  I_3597_S;
wire  I_3599_S;
wire  I_3601_S;
wire  I_3602_D;
wire  I_3602_S;
wire  I_3603_D;
wire  I_3603_G;
wire  I_3603_S;
wire  I_3604_D;
wire  I_3604_S;
wire  I_3605_D;
wire  I_3605_G;
wire  I_3605_S;
wire  I_3606_D;
wire  I_3607_D;
wire  I_3608_D;
wire  I_3609_D;
wire  I_3610_D;
wire  I_3611_D;
wire  I_3612_D;
wire  I_3613_D;
wire  I_3614_D;
wire  I_3615_D;
wire  I_361_G;
wire  I_3621_D;
wire  I_3627_D;
wire  I_362_D;
wire  I_3633_D;
wire  I_3638_D;
wire  I_3638_G;
wire  I_3639_D;
wire  I_3649_D;
wire  I_3649_G;
wire  I_364_D;
wire  I_3651_D;
wire  I_3653_D;
wire  I_3653_S;
wire  I_3655_D;
wire  I_3655_S;
wire  I_3657_D;
wire  I_3658_G;
wire  I_3658_S;
wire  I_3659_G;
wire  I_3659_S;
wire  I_365_D;
wire  I_365_G;
wire  I_3660_D;
wire  I_3663_D;
wire  I_3663_S;
wire  I_3664_G;
wire  I_3664_S;
wire  I_3667_D;
wire  I_3667_S;
wire  I_3669_D;
wire  I_3669_S;
wire  I_366_D;
wire  I_3670_D;
wire  I_3670_G;
wire  I_3670_S;
wire  I_3671_D;
wire  I_3671_G;
wire  I_3671_S;
wire  I_3672_S;
wire  I_3673_S;
wire  I_3675_D;
wire  I_3676_D;
wire  I_3677_D;
wire  I_3678_S;
wire  I_3679_S;
wire  I_367_D;
wire  I_367_G;
wire  I_3681_D;
wire  I_3683_D;
wire  I_368_D;
wire  I_3691_D;
wire  I_3692_D;
wire  I_3695_D;
wire  I_3699_D;
wire  I_369_D;
wire  I_369_G;
wire  I_36_D;
wire  I_3701_D;
wire  I_3703_D;
wire  I_370_D;
wire  I_3718_D;
wire  I_371_D;
wire  I_371_G;
wire  I_3720_D;
wire  I_3724_D;
wire  I_3725_D;
wire  I_3727_G;
wire  I_3728_D;
wire  I_372_D;
wire  I_3731_G;
wire  I_3733_G;
wire  I_3735_G;
wire  I_3736_D;
wire  I_3738_D;
wire  I_373_D;
wire  I_3740_D;
wire  I_3742_D;
wire  I_3744_D;
wire  I_3745_D;
wire  I_3746_D;
wire  I_3747_D;
wire  I_3748_D;
wire  I_3751_S;
wire  I_3752_D;
wire  I_3753_D;
wire  I_3755_D;
wire  I_3755_S;
wire  I_3759_S;
wire  I_375_D;
wire  I_3763_S;
wire  I_3765_S;
wire  I_3766_D;
wire  I_3767_D;
wire  I_3767_G;
wire  I_3768_D;
wire  I_3769_D;
wire  I_3770_D;
wire  I_3771_D;
wire  I_3772_D;
wire  I_3773_D;
wire  I_3774_D;
wire  I_3775_D;
wire  I_3781_D;
wire  I_3788_D;
wire  I_3791_D;
wire  I_3793_D;
wire  I_3795_D;
wire  I_3797_D;
wire  I_379_G;
wire  I_3808_D;
wire  I_3809_D;
wire  I_3810_D;
wire  I_3811_D;
wire  I_3813_D;
wire  I_3813_S;
wire  I_3815_D;
wire  I_3815_S;
wire  I_3816_D;
wire  I_3817_D;
wire  I_3818_D;
wire  I_3819_G;
wire  I_381_G;
wire  I_3820_D;
wire  I_3823_D;
wire  I_3823_S;
wire  I_3824_G;
wire  I_3824_S;
wire  I_3825_D;
wire  I_3825_S;
wire  I_3827_D;
wire  I_3829_D;
wire  I_3829_S;
wire  I_382_D;
wire  I_3830_D;
wire  I_3830_G;
wire  I_3831_D;
wire  I_3832_S;
wire  I_3833_S;
wire  I_3834_D;
wire  I_3835_D;
wire  I_3836_D;
wire  I_3836_G;
wire  I_3837_D;
wire  I_3838_S;
wire  I_3839_S;
wire  I_3845_D;
wire  I_3847_D;
wire  I_3847_G;
wire  I_3850_D;
wire  I_3851_G;
wire  I_3852_D;
wire  I_3854_D;
wire  I_3855_D;
wire  I_3855_G;
wire  I_3856_D;
wire  I_3857_D;
wire  I_3857_G;
wire  I_3859_D;
wire  I_385_D;
wire  I_3861_D;
wire  I_3867_D;
wire  I_3869_D;
wire  I_3872_D;
wire  I_3874_D;
wire  I_387_S;
wire  I_3880_D;
wire  I_3882_D;
wire  I_3883_D;
wire  I_3884_D;
wire  I_3887_D;
wire  I_3889_D;
wire  I_3893_G;
wire  I_3894_D;
wire  I_3896_D;
wire  I_389_S;
wire  I_3902_D;
wire  I_3904_D;
wire  I_3904_S;
wire  I_3905_G;
wire  I_3905_S;
wire  I_3906_D;
wire  I_3906_S;
wire  I_3907_G;
wire  I_3907_S;
wire  I_3908_D;
wire  I_3909_D;
wire  I_390_D;
wire  I_3910_D;
wire  I_3911_D;
wire  I_3911_G;
wire  I_3912_D;
wire  I_3913_S;
wire  I_3915_G;
wire  I_3915_S;
wire  I_3917_S;
wire  I_3919_S;
wire  I_3921_S;
wire  I_3923_G;
wire  I_3923_S;
wire  I_3924_D;
wire  I_3924_S;
wire  I_3925_D;
wire  I_3925_G;
wire  I_3925_S;
wire  I_3926_D;
wire  I_3926_S;
wire  I_3927_G;
wire  I_3927_S;
wire  I_3928_D;
wire  I_3929_D;
wire  I_3930_D;
wire  I_3931_D;
wire  I_3932_D;
wire  I_3933_D;
wire  I_3933_G;
wire  I_3934_D;
wire  I_3935_D;
wire  I_3937_D;
wire  I_3939_D;
wire  I_393_S;
wire  I_394_D;
wire  I_3950_D;
wire  I_3950_G;
wire  I_3953_D;
wire  I_3955_D;
wire  I_3956_D;
wire  I_3956_G;
wire  I_3958_D;
wire  I_3958_G;
wire  I_395_D;
wire  I_3961_D;
wire  I_3968_G;
wire  I_3968_S;
wire  I_3969_S;
wire  I_396_D;
wire  I_396_S;
wire  I_3970_G;
wire  I_3970_S;
wire  I_3971_G;
wire  I_3971_S;
wire  I_3972_D;
wire  I_3973_D;
wire  I_3974_D;
wire  I_3974_G;
wire  I_3975_D;
wire  I_3976_D;
wire  I_3977_D;
wire  I_3977_G;
wire  I_3979_D;
wire  I_397_D;
wire  I_397_G;
wire  I_397_S;
wire  I_3980_D;
wire  I_3980_G;
wire  I_3981_D;
wire  I_3982_G;
wire  I_3983_D;
wire  I_3983_G;
wire  I_3983_S;
wire  I_3985_D;
wire  I_3985_S;
wire  I_3986_G;
wire  I_3986_S;
wire  I_3987_G;
wire  I_3987_S;
wire  I_3988_G;
wire  I_3988_S;
wire  I_3989_G;
wire  I_3989_S;
wire  I_398_D;
wire  I_398_S;
wire  I_3990_G;
wire  I_3990_S;
wire  I_3991_G;
wire  I_3991_S;
wire  I_3992_G;
wire  I_3992_S;
wire  I_3993_G;
wire  I_3993_S;
wire  I_3994_D;
wire  I_3995_D;
wire  I_3996_D;
wire  I_3997_D;
wire  I_3999_D;
wire  I_3999_G;
wire  I_399_D;
wire  I_399_G;
wire  I_399_S;
wire  I_3_D;
wire  I_3_G;
wire  I_400_D;
wire  I_400_S;
wire  I_401_D;
wire  I_401_G;
wire  I_401_S;
wire  I_402_D;
wire  I_402_S;
wire  I_403_D;
wire  I_403_G;
wire  I_403_S;
wire  I_404_S;
wire  I_405_G;
wire  I_405_S;
wire  I_409_S;
wire  I_40_D;
wire  I_410_D;
wire  I_410_S;
wire  I_411_D;
wire  I_411_G;
wire  I_411_S;
wire  I_415_S;
wire  I_418_D;
wire  I_418_G;
wire  I_419_D;
wire  I_41_D;
wire  I_41_G;
wire  I_421_D;
wire  I_423_D;
wire  I_426_D;
wire  I_426_G;
wire  I_429_D;
wire  I_42_D;
wire  I_430_D;
wire  I_430_G;
wire  I_431_D;
wire  I_432_D;
wire  I_432_G;
wire  I_433_D;
wire  I_434_D;
wire  I_434_G;
wire  I_435_D;
wire  I_437_D;
wire  I_439_D;
wire  I_43_D;
wire  I_43_G;
wire  I_443_D;
wire  I_445_D;
wire  I_447_D;
wire  I_448_D;
wire  I_449_D;
wire  I_44_D;
wire  I_450_D;
wire  I_450_G;
wire  I_450_S;
wire  I_451_D;
wire  I_451_G;
wire  I_451_S;
wire  I_453_D;
wire  I_453_S;
wire  I_455_D;
wire  I_456_D;
wire  I_457_D;
wire  I_458_S;
wire  I_459_G;
wire  I_459_S;
wire  I_45_D;
wire  I_45_G;
wire  I_460_G;
wire  I_460_S;
wire  I_461_S;
wire  I_462_D;
wire  I_462_G;
wire  I_462_S;
wire  I_463_D;
wire  I_463_G;
wire  I_463_S;
wire  I_464_D;
wire  I_464_G;
wire  I_464_S;
wire  I_465_D;
wire  I_465_G;
wire  I_465_S;
wire  I_466_D;
wire  I_466_G;
wire  I_466_S;
wire  I_467_D;
wire  I_467_G;
wire  I_467_S;
wire  I_468_D;
wire  I_469_D;
wire  I_46_D;
wire  I_471_D;
wire  I_471_S;
wire  I_473_D;
wire  I_475_D;
wire  I_477_D;
wire  I_477_S;
wire  I_479_D;
wire  I_47_D;
wire  I_47_G;
wire  I_482_D;
wire  I_483_D;
wire  I_483_G;
wire  I_48_D;
wire  I_493_G;
wire  I_494_D;
wire  I_495_D;
wire  I_495_G;
wire  I_496_D;
wire  I_497_D;
wire  I_497_G;
wire  I_498_D;
wire  I_499_D;
wire  I_499_G;
wire  I_49_D;
wire  I_49_G;
wire  I_500_D;
wire  I_501_D;
wire  I_501_G;
wire  I_503_D;
wire  I_503_G;
wire  I_505_D;
wire  I_507_G;
wire  I_509_D;
wire  I_50_D;
wire  I_511_D;
wire  I_513_D;
wire  I_516_D;
wire  I_51_D;
wire  I_51_G;
wire  I_520_D;
wire  I_522_D;
wire  I_524_D;
wire  I_525_D;
wire  I_526_D;
wire  I_527_D;
wire  I_527_G;
wire  I_528_D;
wire  I_529_D;
wire  I_529_G;
wire  I_52_D;
wire  I_530_D;
wire  I_531_D;
wire  I_531_G;
wire  I_532_D;
wire  I_533_D;
wire  I_533_G;
wire  I_535_G;
wire  I_539_G;
wire  I_53_D;
wire  I_53_G;
wire  I_543_G;
wire  I_544_D;
wire  I_545_D;
wire  I_546_D;
wire  I_547_D;
wire  I_549_S;
wire  I_550_D;
wire  I_552_D;
wire  I_553_D;
wire  I_554_D;
wire  I_555_D;
wire  I_556_S;
wire  I_557_G;
wire  I_557_S;
wire  I_558_D;
wire  I_558_S;
wire  I_559_D;
wire  I_559_G;
wire  I_559_S;
wire  I_55_G;
wire  I_560_D;
wire  I_560_S;
wire  I_561_D;
wire  I_561_G;
wire  I_561_S;
wire  I_562_D;
wire  I_562_S;
wire  I_563_D;
wire  I_563_G;
wire  I_563_S;
wire  I_564_D;
wire  I_564_S;
wire  I_565_D;
wire  I_565_G;
wire  I_565_S;
wire  I_566_D;
wire  I_566_S;
wire  I_567_D;
wire  I_567_G;
wire  I_567_S;
wire  I_56_D;
wire  I_571_G;
wire  I_572_D;
wire  I_573_D;
wire  I_575_S;
wire  I_57_D;
wire  I_57_G;
wire  I_581_D;
wire  I_583_D;
wire  I_584_D;
wire  I_584_G;
wire  I_586_D;
wire  I_586_G;
wire  I_588_D;
wire  I_588_G;
wire  I_589_D;
wire  I_590_D;
wire  I_590_G;
wire  I_591_D;
wire  I_592_D;
wire  I_592_G;
wire  I_593_D;
wire  I_594_D;
wire  I_594_G;
wire  I_595_D;
wire  I_596_D;
wire  I_596_G;
wire  I_597_D;
wire  I_59_D;
wire  I_601_D;
wire  I_603_D;
wire  I_607_D;
wire  I_608_D;
wire  I_609_D;
wire  I_610_D;
wire  I_611_D;
wire  I_613_D;
wire  I_613_S;
wire  I_615_D;
wire  I_616_S;
wire  I_617_G;
wire  I_617_S;
wire  I_618_S;
wire  I_619_G;
wire  I_619_S;
wire  I_620_D;
wire  I_620_G;
wire  I_620_S;
wire  I_621_D;
wire  I_621_G;
wire  I_621_S;
wire  I_622_D;
wire  I_622_G;
wire  I_622_S;
wire  I_623_D;
wire  I_623_G;
wire  I_623_S;
wire  I_624_D;
wire  I_624_G;
wire  I_624_S;
wire  I_625_D;
wire  I_625_G;
wire  I_625_S;
wire  I_626_D;
wire  I_626_G;
wire  I_626_S;
wire  I_627_D;
wire  I_627_G;
wire  I_627_S;
wire  I_628_D;
wire  I_628_G;
wire  I_628_S;
wire  I_629_D;
wire  I_629_G;
wire  I_629_S;
wire  I_631_D;
wire  I_633_D;
wire  I_634_D;
wire  I_635_D;
wire  I_637_D;
wire  I_638_G;
wire  I_638_S;
wire  I_639_S;
wire  I_640_D;
wire  I_641_D;
wire  I_641_G;
wire  I_648_D;
wire  I_649_D;
wire  I_649_G;
wire  I_652_D;
wire  I_653_D;
wire  I_653_G;
wire  I_654_D;
wire  I_655_D;
wire  I_655_G;
wire  I_656_D;
wire  I_657_D;
wire  I_657_G;
wire  I_658_D;
wire  I_659_D;
wire  I_659_G;
wire  I_65_S;
wire  I_660_D;
wire  I_661_D;
wire  I_661_G;
wire  I_667_D;
wire  I_670_D;
wire  I_671_D;
wire  I_671_G;
wire  I_674_D;
wire  I_675_D;
wire  I_676_D;
wire  I_67_D;
wire  I_67_S;
wire  I_680_D;
wire  I_681_D;
wire  I_681_G;
wire  I_682_D;
wire  I_684_D;
wire  I_685_D;
wire  I_685_G;
wire  I_686_D;
wire  I_687_D;
wire  I_687_G;
wire  I_688_D;
wire  I_689_D;
wire  I_689_G;
wire  I_690_D;
wire  I_691_D;
wire  I_691_G;
wire  I_692_D;
wire  I_693_D;
wire  I_693_G;
wire  I_698_D;
wire  I_699_D;
wire  I_69_S;
wire  I_700_D;
wire  I_705_D;
wire  I_707_S;
wire  I_709_S;
wire  I_70_D;
wire  I_710_D;
wire  I_713_S;
wire  I_714_D;
wire  I_715_D;
wire  I_716_D;
wire  I_716_S;
wire  I_717_D;
wire  I_717_G;
wire  I_717_S;
wire  I_718_D;
wire  I_718_S;
wire  I_719_D;
wire  I_719_G;
wire  I_719_S;
wire  I_720_D;
wire  I_720_S;
wire  I_721_D;
wire  I_721_G;
wire  I_721_S;
wire  I_722_D;
wire  I_722_S;
wire  I_723_D;
wire  I_723_G;
wire  I_723_S;
wire  I_727_D;
wire  I_729_S;
wire  I_72_D;
wire  I_72_S;
wire  I_730_S;
wire  I_731_G;
wire  I_731_S;
wire  I_733_S;
wire  I_735_D;
wire  I_738_D;
wire  I_738_G;
wire  I_739_D;
wire  I_73_D;
wire  I_73_G;
wire  I_73_S;
wire  I_741_D;
wire  I_743_D;
wire  I_747_D;
wire  I_748_D;
wire  I_748_G;
wire  I_749_D;
wire  I_74_D;
wire  I_74_S;
wire  I_750_D;
wire  I_750_G;
wire  I_751_D;
wire  I_752_D;
wire  I_752_G;
wire  I_753_D;
wire  I_754_D;
wire  I_754_G;
wire  I_755_D;
wire  I_759_D;
wire  I_75_D;
wire  I_75_G;
wire  I_75_S;
wire  I_763_D;
wire  I_765_D;
wire  I_767_D;
wire  I_768_D;
wire  I_769_D;
wire  I_76_D;
wire  I_76_S;
wire  I_770_D;
wire  I_770_G;
wire  I_770_S;
wire  I_771_D;
wire  I_771_G;
wire  I_771_S;
wire  I_773_D;
wire  I_773_S;
wire  I_775_D;
wire  I_777_D;
wire  I_778_G;
wire  I_778_S;
wire  I_779_S;
wire  I_77_D;
wire  I_77_G;
wire  I_77_S;
wire  I_780_D;
wire  I_780_G;
wire  I_780_S;
wire  I_781_D;
wire  I_781_G;
wire  I_781_S;
wire  I_782_D;
wire  I_782_G;
wire  I_782_S;
wire  I_783_D;
wire  I_783_G;
wire  I_783_S;
wire  I_784_D;
wire  I_784_G;
wire  I_784_S;
wire  I_785_D;
wire  I_785_G;
wire  I_785_S;
wire  I_786_D;
wire  I_786_G;
wire  I_786_S;
wire  I_787_D;
wire  I_787_G;
wire  I_787_S;
wire  I_789_D;
wire  I_78_D;
wire  I_78_S;
wire  I_791_D;
wire  I_793_D;
wire  I_795_D;
wire  I_797_D;
wire  I_798_G;
wire  I_798_S;
wire  I_799_S;
wire  I_79_D;
wire  I_79_G;
wire  I_79_S;
wire  I_802_D;
wire  I_803_D;
wire  I_803_G;
wire  I_809_D;
wire  I_80_D;
wire  I_80_S;
wire  I_810_D;
wire  I_811_D;
wire  I_811_G;
wire  I_812_D;
wire  I_813_D;
wire  I_813_G;
wire  I_814_D;
wire  I_815_D;
wire  I_815_G;
wire  I_816_D;
wire  I_817_D;
wire  I_817_G;
wire  I_818_D;
wire  I_819_D;
wire  I_819_G;
wire  I_81_D;
wire  I_81_G;
wire  I_81_S;
wire  I_821_D;
wire  I_825_D;
wire  I_827_D;
wire  I_82_D;
wire  I_82_S;
wire  I_833_D;
wire  I_836_D;
wire  I_83_D;
wire  I_83_G;
wire  I_83_S;
wire  I_842_D;
wire  I_843_D;
wire  I_843_G;
wire  I_844_D;
wire  I_845_D;
wire  I_845_G;
wire  I_846_D;
wire  I_847_D;
wire  I_847_G;
wire  I_848_D;
wire  I_849_D;
wire  I_849_G;
wire  I_850_D;
wire  I_851_D;
wire  I_851_G;
wire  I_852_D;
wire  I_853_D;
wire  I_855_D;
wire  I_858_D;
wire  I_859_D;
wire  I_85_G;
wire  I_861_G;
wire  I_862_D;
wire  I_864_D;
wire  I_865_D;
wire  I_866_D;
wire  I_867_D;
wire  I_869_S;
wire  I_870_D;
wire  I_873_D;
wire  I_874_D;
wire  I_874_S;
wire  I_875_D;
wire  I_875_G;
wire  I_875_S;
wire  I_876_D;
wire  I_876_S;
wire  I_877_D;
wire  I_877_G;
wire  I_877_S;
wire  I_878_D;
wire  I_878_S;
wire  I_879_D;
wire  I_879_G;
wire  I_879_S;
wire  I_87_G;
wire  I_880_D;
wire  I_880_S;
wire  I_881_D;
wire  I_881_G;
wire  I_881_S;
wire  I_882_D;
wire  I_882_S;
wire  I_883_D;
wire  I_883_G;
wire  I_883_S;
wire  I_884_S;
wire  I_885_G;
wire  I_885_S;
wire  I_88_D;
wire  I_88_S;
wire  I_890_S;
wire  I_891_G;
wire  I_891_S;
wire  I_894_D;
wire  I_89_D;
wire  I_89_G;
wire  I_89_S;
wire  I_8_D;
wire  I_901_D;
wire  I_903_D;
wire  I_906_D;
wire  I_906_G;
wire  I_907_D;
wire  I_908_D;
wire  I_908_G;
wire  I_909_D;
wire  I_910_D;
wire  I_910_G;
wire  I_911_D;
wire  I_912_D;
wire  I_912_G;
wire  I_913_D;
wire  I_914_D;
wire  I_914_G;
wire  I_915_D;
wire  I_917_D;
wire  I_919_D;
wire  I_91_G;
wire  I_921_D;
wire  I_923_D;
wire  I_925_D;
wire  I_928_D;
wire  I_929_D;
wire  I_930_D;
wire  I_931_D;
wire  I_933_D;
wire  I_933_S;
wire  I_935_D;
wire  I_937_D;
wire  I_938_D;
wire  I_938_G;
wire  I_938_S;
wire  I_939_D;
wire  I_939_G;
wire  I_939_S;
wire  I_93_S;
wire  I_940_D;
wire  I_940_G;
wire  I_940_S;
wire  I_941_D;
wire  I_941_G;
wire  I_941_S;
wire  I_942_D;
wire  I_942_G;
wire  I_942_S;
wire  I_943_D;
wire  I_943_G;
wire  I_943_S;
wire  I_944_D;
wire  I_944_G;
wire  I_944_S;
wire  I_945_D;
wire  I_945_G;
wire  I_945_S;
wire  I_946_D;
wire  I_946_G;
wire  I_946_S;
wire  I_947_D;
wire  I_947_G;
wire  I_947_S;
wire  I_948_D;
wire  I_949_D;
wire  I_951_D;
wire  I_953_D;
wire  I_954_D;
wire  I_955_D;
wire  I_957_D;
wire  I_957_S;
wire  I_959_D;
wire  I_95_D;
wire  I_95_G;
wire  I_960_D;
wire  I_961_D;
wire  I_961_G;
wire  I_969_D;
wire  I_970_D;
wire  I_971_D;
wire  I_971_G;
wire  I_972_D;
wire  I_973_D;
wire  I_973_G;
wire  I_975_D;
wire  I_976_D;
wire  I_977_D;
wire  I_977_G;
wire  I_978_D;
wire  I_979_D;
wire  I_979_G;
wire  I_983_D;
wire  I_989_D;
wire  I_994_D;
wire  I_995_D;
wire  I_998_D;
wire  I_99_D;
wire  I_9_D;
wire  I_9_G;

	nand auto_290(I_33_D, I_3_G, I_65_S);
	not auto_291(I_1033_D, I_969_D); // NMOS strength = 2
	nand auto_292(I_1039_D, I_1741_S, I_1997_D);
	not auto_293(I_1045_D, I_983_D); // NMOS strength = 3
	not auto_294(I_1401_D, I_953_D); // NMOS strength = 2
	not auto_295(I_1397_D, I_925_D); // NMOS strength = 2
	nand auto_296(I_1087_D, I_1117_D, I_959_D);
	not auto_297(I_1025_D, I_1025_G); // NMOS strength = 2
	not auto_298(I_1027_S, I_1249_D);
	nand auto_299(I_1029_D, I_1093_D, I_1187_S);
	not auto_300(I_1093_S, I_1095_D);
	not auto_301(I_1049_S, I_1401_D);
	not auto_302(I_1051_S, I_445_D); // NMOS strength = 2
	not auto_303(I_1055_S, I_1087_D);
	nand auto_304(I_1089_D, I_1667_D, I_1153_G);
	nand auto_305(I_1091_D, I_389_S, I_1985_S);
	nand auto_306(I_1103_D, I_975_D, I_2471_S);
	nand auto_307(I_1115_D, I_1275_D, I_1205_D);
	not auto_308(I_1097_S, I_715_D);
	not auto_309(I_1099_S, I_1258_G);
	not auto_310(I_1101_S, I_1973_D);
	nand auto_311(I_1113_S, I_1529_D, I_1529_D);
	not auto_312(I_1187_S, I_1539_D); // NMOS strength = 3
	not auto_313(I_1221_D, I_1189_D);
	nand auto_314(I_1223_D, I_1187_S, I_1253_S);
	not auto_315(I_1225_D, I_1259_S);
	not auto_316(I_1227_D, I_1195_D);
	nand auto_317(I_2071_S, I_1103_D, I_1039_D);
	not auto_318(I_1139_D, I_1269_S);
	not auto_319(I_1237_D, I_1205_D);
	not auto_320(I_1239_D, I_1207_D);
	nand auto_321(I_1211_D, I_1051_S, I_735_D, I_1397_D);
	nand auto_322(I_1213_D, I_957_S, I_511_D, I_477_S);
	not auto_323(I_1279_S, I_1119_D);
	nand auto_324(I_1185_D, I_1153_G, I_1185_G);
	nand auto_325(I_1189_D, I_1187_S, I_1253_D);
	not auto_326(I_1259_S, I_1193_G); // NMOS strength = 2
	not auto_327(I_1195_D, I_1259_D); // NMOS strength = 2
	not auto_328(I_1269_S, I_1267_D); // NMOS strength = 2
	not auto_329(I_1205_D, I_1269_D); // NMOS strength = 2
	not auto_330(I_1207_D, I_1271_D); // NMOS strength = 2
	not auto_331(I_151_D, I_151_G);
	not auto_332(I_1253_S, I_1255_D);
	nand auto_333(I_1209_S, I_1435_D, I_1435_D);
	not auto_334(I_1247_D, I_1279_S);
	not auto_335(I_1249_D, I_1251_D); // NMOS strength = 2
	nand auto_336(I_1251_D, I_1091_D, I_1250_G);
	not auto_337(I_1417_S, I_1260_G);
	not auto_338(I_1267_S, I_1262_G);
	nand auto_339(I_1275_D, I_1307_D, I_735_D);
	not auto_340(I_1407_D, I_1343_D);
	nand auto_341(I_1273_S, I_1209_S, I_1209_S);
	not auto_342(I_1283_D, I_1345_D);
	not auto_343(I_1381_D, I_1349_D);
	nand auto_344(I_1383_D, I_1187_S, I_1413_S);
	not auto_345(I_1385_D, I_1419_S);
	not auto_346(I_1387_D, I_1355_D);
	not auto_347(I_1295_D, I_1997_D);
	not auto_348(I_1297_D, I_1999_D);
	not auto_349(I_1301_D, I_735_D);
	not auto_350(I_1335_D, I_1431_D); // NMOS strength = 2
	not auto_351(I_1307_D, I_957_S);
	nand auto_352(I_1309_D, I_1369_S, I_1369_S);
	not auto_353(I_131_S, I_67_S);
	nand auto_354(I_1343_D, I_1311_G, I_1439_D);
	nand auto_355(I_1345_D, I_1313_G, I_1409_D);
	not auto_356(I_1347_D, I_1345_D); // NMOS strength = 2
	nand auto_357(I_1349_D, I_1187_S, I_1413_D);
	not auto_358(I_1419_S, I_1417_D); // NMOS strength = 2
	not auto_359(I_1355_D, I_1419_D); // NMOS strength = 2
	nand auto_360(I_1359_D, I_3111_S, I_1997_D);
	nand auto_361(I_1331_D, I_1365_S, I_1365_S);
	not auto_362(I_1413_S, I_1415_D);
	not auto_363(I_1361_S, I_2071_S);
	nand auto_364(I_1365_S, I_1523_S, I_1523_S);
	not auto_365(I_1399_D, I_1335_D);
	nand auto_366(I_1369_S, I_1273_S, I_1273_S);
	not auto_367(I_1373_S, I_1247_D);
	nand auto_368(I_1409_D, I_1409_G, I_1408_G);
	not auto_369(I_1420_S, I_1101_S);
	nand auto_370(I_1423_D, I_1295_D, I_2631_S);
	nor auto_371(I_1435_D, I_1307_D, I_1373_S, I_1051_S);
	not auto_372(I_1411_S, I_1671_S);
	nor auto_373(I_1913_S, I_1397_D, I_735_D);
	not auto_374(I_1537_D, I_1571_S);
	not auto_375(I_1539_D, I_1507_D);
	not auto_376(I_1541_D, I_1575_S);
	nand auto_377(I_1573_S, I_1511_S, I_1347_D);
	nand auto_378(I_1483_D, I_1195_D, VDD);
	nand auto_379(I_1518_D, I_1359_D, I_1423_D);
	not auto_380(I_1491_D, I_1427_D); // NMOS strength = 2
	not auto_381(I_1461_D, I_1525_D);
	not auto_382(I_1559_D, I_1593_S);
	not auto_383(I_1561_D, I_1529_D);
	nand auto_384(I_1499_D, I_1997_D, I_1051_S);
	not auto_385(I_1469_D, I_1213_D);
	nand auto_386(I_1535_D, I_3667_D, I_1758_S, I_1598_S);
	not auto_387(I_1571_S, I_1569_D); // NMOS strength = 2
	not auto_388(I_1507_D, I_1571_D); // NMOS strength = 2
	nand auto_389(I_1575_S, I_1347_D, I_1573_D);
	not auto_390(I_1525_D, I_1429_D); // NMOS strength = 2
	not auto_391(I_1593_S, I_1591_D); // NMOS strength = 2
	not auto_392(I_1529_D, I_1593_D); // NMOS strength = 2
	not auto_393(I_1597_D, I_1627_D); // NMOS strength = 4
	not auto_394(I_1511_S, I_1575_D);
	not auto_395(I_1515_S, I_1483_D);
	not auto_396(I_1523_S, I_1491_D);
	not auto_397(I_1531_S, I_1499_D);
	not auto_398(I_1576_S, I_1051_S);
	nand auto_399(I_1585_D, I_1679_D, I_1518_D);
	not auto_400(I_1588_S, I_1685_D);
	not auto_401(I_1627_D, I_1531_S); // NMOS strength = 3
	not auto_402(I_1598_S, I_1597_D);
	not auto_403(I_1589_S, I_1588_S);
	not auto_404(I_1599_S, I_1598_S);
	not auto_405(I_1697_D, I_1731_S);
	not auto_406(I_1699_D, I_1667_D);
	not auto_407(I_1701_D, I_1735_S);
	nand auto_408(I_1733_S, I_1347_D, I_1671_S);
	not auto_409(I_1609_D, I_1249_D);
	nor auto_410(I_1648_D, I_1518_D, I_1679_D);
	not auto_411(I_1623_D, I_1687_S);
	not auto_412(I_1689_D, I_1879_D); // NMOS strength = 3
	nand auto_413(I_1693_D, I_1535_D, I_1695_D, I_1855_D);
	nand auto_414(I_1695_D, I_1598_S, I_1631_G, I_1759_S);
	not auto_415(I_1731_S, I_1729_D); // NMOS strength = 2
	not auto_416(I_1667_D, I_1731_D); // NMOS strength = 2
	nand auto_417(I_1735_S, I_1347_D, I_1733_D);
	nand auto_418(I_1673_D, I_1515_S, I_1249_D);
	nand auto_419(I_1679_D, I_1807_D, I_1743_D);
	nand auto_420(I_261_D, I_1187_S, I_229_S);
	not auto_421(I_1685_D, I_151_D);
	not auto_422(I_1755_D, I_1627_D); // NMOS strength = 4
	not auto_423(I_263_D, I_293_S);
	not auto_424(I_1671_S, I_1735_D);
	not auto_425(I_1681_S, I_1648_D);
	not auto_426(I_1687_S, I_1685_D);
	nand auto_427(I_1737_D, I_1515_S, I_1609_D);
	nand auto_428(I_235_D, I_458_S, I_297_S, I_618_S);
	nand auto_429(I_1743_D, I_1839_S, I_1741_S);
	not auto_430(I_1748_S, I_1751_S);
	not auto_431(I_1750_S, I_151_D);
	not auto_432(I_1752_S, I_1751_S);
	not auto_433(I_1757_D, I_1915_S); // NMOS strength = 2
	not auto_434(I_1758_S, I_1821_D);
	not auto_435(I_1741_S, I_3013_S);
	not auto_436(I_1749_S, I_1748_S);
	not auto_437(I_1751_S, I_1750_S);
	not auto_438(I_1753_S, I_1752_S);
	not auto_439(I_1759_S, I_1758_S);
	not auto_440(I_1761_D, I_1761_G);
	not auto_441(I_1763_D, I_1831_S);
	not auto_442(I_1861_D, I_1895_S);
	nand auto_443(I_1893_S, I_1347_D, I_1831_S);
	nand auto_444(I_1832_D, I_1737_D, I_1673_D);
	nand auto_445(I_1807_D, I_3431_S, I_2253_D);
	nand auto_446(I_2065_S, I_1585_D, I_1681_S);
	nand auto_447(I_1845_D, I_1051_S, I_1397_D, I_457_D);
	not auto_448(I_1879_D, I_1847_D);
	not auto_449(I_1881_D, I_1911_S);
	not auto_450(I_1821_D, I_1853_S); // NMOS strength = 4
	nand auto_451(I_1855_D, I_1758_S, I_1599_S, I_1901_D);
	not auto_452(I_1825_D, I_1345_D); // NMOS strength = 2
	nand auto_453(I_1891_S, I_1763_D, I_2311_S, I_1923_D, I_2151_S);
	nand auto_454(I_1895_S, I_1347_D, I_1893_D);
	not auto_455(I_245_D, I_277_D); // NMOS strength = 3
	not auto_456(I_1847_D, I_1911_D); // NMOS strength = 2
	not auto_457(I_1911_S, I_1913_D); // NMOS strength = 2
	not auto_458(I_279_D, I_247_D);
	not auto_459(I_1831_S, I_1895_D);
	not auto_460(I_1839_S, I_2253_D);
	not auto_461(I_2033_D, I_2065_S);
	not auto_462(I_1843_S, I_1425_S);
	not auto_463(I_185_D, I_281_D);
	not auto_464(I_1853_S, I_1279_S); // NMOS strength = 2
	nand auto_465(I_1889_D, I_1987_D, I_1888_G);
	nand auto_466(I_1901_D, I_2157_S, I_101_D);
	not auto_467(I_251_S, I_347_D); // NMOS strength = 3
	not auto_468(I_1906_S, I_1843_S);
	not auto_469(I_1908_S, I_503_D);
	nand auto_470(I_1917_D, I_1693_D, I_1949_D);
	not auto_471(I_1919_D, I_2077_D); // NMOS strength = 2
	nand auto_472(I_285_D, I_159_S, I_157_D);
	nor auto_473(I_1899_S, I_873_D, I_101_D);
	nor auto_474(I_1915_S, I_1879_D, I_1853_S);
	nand auto_475(I_2209_S, I_1985_S, I_1921_G);
	not auto_476(I_1923_D, I_1991_S);
	not auto_477(I_2021_D, I_2055_S);
	nand auto_478(I_2053_S, I_1347_D, I_1991_S);
	nand auto_479(I_225_D, auto_net_1, I_289_D);
	or auto_480(auto_net_1, I_1832_D, I_227_D);
	nor auto_481(I_1962_D, I_1899_S, auto_net_2);
	and auto_482(auto_net_2, I_101_D, I_873_D);
	not auto_483(I_1997_D, I_2317_S); // NMOS strength = 3
	not auto_484(I_1973_D, I_1943_D); // NMOS strength = 2
	not auto_485(I_1943_D, I_1309_D);
	not auto_486(I_2009_D, I_1879_D); // NMOS strength = 3
	not auto_487(I_1949_D, I_1689_D);
	nand auto_488(I_227_D, I_355_D, I_291_D);
	nand auto_489(I_2015_D, I_2238_S, I_3669_D, I_2078_S);
	nand auto_490(I_1987_D, I_2115_D, I_2051_D);
	nand auto_491(I_2055_S, I_1347_D, I_2053_D);
	not auto_492(I_1969_D, I_1906_S);
	not auto_493(I_2007_D, I_1973_D); // NMOS strength = 2
	nand auto_494(I_2011_D, I_2139_D, I_2075_D);
	nand auto_495(I_2013_D, I_1689_D, I_2011_D);
	not auto_496(I_1985_S, I_2049_D);
	nand auto_497(I_293_S, I_1187_S, I_295_D);
	not auto_498(I_1991_S, I_2055_D);
	not auto_499(I_2001_S, I_1969_D);
	nand auto_500(I_2051_D, I_2050_G, I_2147_S);
	not auto_501(I_2058_S, I_2699_D);
	nand auto_502(I_2063_D, I_2159_S, I_2062_G);
	nand auto_503(I_2069_D, I_2133_G, I_1518_D);
	nand auto_504(I_2075_D, I_2171_S, I_2071_D);
	nand auto_505(I_2077_D, I_1917_D, I_2013_D);
	not auto_506(I_2078_S, I_1597_D);
	not auto_507(I_2079_S, I_2078_S);
	nand auto_508(I_2113_D, I_2209_D, I_2113_G);
	nand auto_509(I_2115_D, I_2083_G, I_1033_D);
	not auto_510(I_2181_D, I_2215_S);
	nand auto_511(I_2213_S, I_2151_S, I_1347_D);
	nor auto_512(I_2154_D, I_3562_D, I_2539_S, I_2058_S);
	nand auto_513(I_2127_D, I_3271_S, I_1997_D);
	nor auto_514(I_2132_D, I_1518_D, I_2133_G);
	not auto_515(I_2103_D, I_2231_D);
	not auto_516(I_2105_D, I_2073_D);
	nand auto_517(I_2139_D, I_2169_D, I_1755_D);
	nand auto_518(I_2173_D, I_2015_D, I_2175_D, I_2335_D);
	nand auto_519(I_2175_D, I_2078_S, I_3923_S, I_2239_S);
	nand auto_520(I_2215_S, I_2213_D, I_1347_D);
	not auto_521(I_2169_D, I_2105_D); // NMOS strength = 2
	not auto_522(I_2177_D, I_2113_D);
	not auto_523(I_2147_S, I_1033_D);
	not auto_524(I_247_D, I_311_D); // NMOS strength = 2
	not auto_525(I_2151_S, I_2215_D);
	not auto_526(I_2157_S, I_873_D);
	not auto_527(I_2159_S, I_1997_D);
	not auto_528(I_2165_S, I_2132_D);
	not auto_529(I_2167_S, I_2071_S);
	not auto_530(I_281_D, I_153_D); // NMOS strength = 2
	not auto_531(I_2171_S, I_1755_D);
	nand auto_532(I_2211_D, I_2213_S, I_2053_S);
	not auto_533(I_2253_D, I_2317_S); // NMOS strength = 3
	nand auto_534(I_2225_D, I_1999_D, I_2319_D);
	nand auto_535(I_2235_D, I_2267_D, I_2549_D);
	nand auto_536(I_2237_D, I_2269_D, I_2173_D);
	not auto_537(I_2238_S, I_1821_D);
	not auto_538(I_2219_S, I_2154_D);
	not auto_539(I_2239_S, I_2238_S);
	nand auto_540(I_2529_S, I_2305_S, I_2241_G);
	nand auto_541(I_2275_D, I_2311_S, I_2211_D);
	not auto_542(I_2341_D, I_2375_S);
	nand auto_543(I_2373_S, I_2311_S, I_1347_D);
	nor auto_544(I_2288_D, I_1999_D, I_2319_D);
	nand auto_545(I_2549_S, I_2165_S, I_2069_D);
	not auto_546(I_2263_D, I_2231_S);
	not auto_547(I_2265_D, I_2233_D);
	not auto_548(I_2267_D, I_1755_D);
	not auto_549(I_2269_D, I_2009_D);
	nand auto_550(I_2335_D, I_2079_S, I_2238_S, VDD);
	nand auto_551(I_2375_S, I_1347_D, I_2373_D);
	nand auto_552(I_2319_D, I_2383_D, I_2447_D);
	not auto_553(I_229_S, I_293_D);
	not auto_554(I_2329_D, I_2265_D); // NMOS strength = 2
	nand auto_555(I_2331_D, I_1755_D, I_2329_D);
	not auto_556(I_2521_D, I_23_G);
	nand auto_557(I_2333_D, I_2395_D, I_2009_D);
	not auto_558(I_2305_S, I_2369_D);
	not auto_559(I_2311_S, I_2375_D);
	not auto_560(I_2317_S, I_3499_D);
	not auto_561(I_2321_S, I_2288_D);
	not auto_562(I_2517_D, I_2549_S);
	not auto_563(I_2389_S, I_2263_D);
	nand auto_564(I_2383_D, I_3111_S, I_2479_S);
	nand auto_565(I_2391_D, I_1265_D, I_2311_S);
	nand auto_566(I_2395_D, I_2331_D, I_2235_D);
	nand auto_567(I_2397_D, I_2237_D, I_2333_D);
	not auto_568(I_2399_D, I_2397_D); // NMOS strength = 2
	nor auto_569(I_2371_S, I_2632_D, I_2370_G);
	nor auto_570(I_2379_S, I_3499_D, I_3337_D);
	nand auto_571(I_2433_D, I_2529_D, I_2433_G);
	not auto_572(I_2501_D, I_2535_S);
	nand auto_573(I_2533_S, I_3241_D, I_2471_S);
	nand auto_574(I_2447_D, I_3337_D, I_2253_D);
	nand auto_575(I_2705_S, I_2225_D, I_2321_S);
	nor auto_576(I_2454_D, I_2311_S, I_1265_D);
	not auto_577(I_2425_D, I_2393_D);
	not auto_578(I_2427_D, I_1755_D);
	not auto_579(I_2429_D, I_2009_D);
	nand auto_580(I_2495_D, I_3036_S, I_2718_S, I_2558_S);
	nand auto_581(I_2535_S, I_3241_D, I_2533_D);
	not auto_582(I_2453_D, I_2389_S);
	not auto_583(I_2489_D, I_2425_D); // NMOS strength = 2
	nand auto_584(I_2491_D, I_1755_D, I_2489_D);
	nand auto_585(I_2493_D, I_2009_D, I_2650_D);
	not auto_586(I_2497_D, I_2433_D);
	not auto_587(I_2471_S, I_2535_D);
	not auto_588(I_2479_S, I_2253_D);
	not auto_589(I_2673_D, I_2705_S);
	not auto_590(I_2485_S, I_2453_D);
	not auto_591(I_2487_S, I_2454_D);
	not auto_592(I_2530_S, I_2535_G);
	nand auto_593(I_2555_D, I_2427_D, I_2871_D);
	nand auto_594(I_2557_D, I_2653_D, I_2429_D);
	not auto_595(I_2558_S, I_1597_D);
	not auto_596(I_253_S, I_285_D);
	nor auto_597(I_2539_S, I_3751_S, I_3591_S);
	not auto_598(I_2559_S, I_2558_S);
	nand auto_599(I_2657_D, I_2561_G, I_2625_S);
	not auto_600(I_2661_D, I_2695_S);
	nand auto_601(I_2693_S, I_3241_D, I_2631_S);
	nor auto_602(I_2632_D, I_3653_S, I_3493_S, I_3333_S);
	nand auto_603(I_289_D, I_1832_D, I_227_D);
	nor auto_604(I_2634_D, I_3493_S, I_3751_S, I_3653_S);
	nand auto_605(I_2871_S, I_2487_S, I_2391_D);
	not auto_606(I_2585_D, I_2553_D);
	nand auto_607(I_2650_D, I_2491_D, I_2555_D);
	nand auto_608(I_2653_D, I_2495_D, I_2655_D, I_2815_D);
	nand auto_609(I_291_D, I_387_S, I_549_S);
	nand auto_610(I_2655_D, I_3593_S, I_2558_S, I_2719_S);
	nand auto_611(I_2695_S, I_3241_D, I_2693_D);
	not auto_612(I_2609_D, I_2545_S);
	not auto_613(I_2649_D, I_2585_D); // NMOS strength = 2
	not auto_614(I_2625_S, I_2689_D);
	not auto_615(I_2631_S, I_2695_D);
	not auto_616(I_2641_S, I_2609_D);
	not auto_617(I_2839_D, I_2871_S);
	nand auto_618(I_2699_D, I_2634_D, I_2794_D);
	nand auto_619(I_2715_D, I_2747_D, I_2709_D);
	nand auto_620(I_2717_D, I_2557_D, I_2493_D);
	not auto_621(I_2718_S, I_1821_D);
	not auto_622(I_59_D, I_1115_D); // NMOS strength = 2
	not auto_623(I_2719_S, I_2718_S);
	nand auto_624(I_2753_D, I_2849_D, I_2753_G);
	not auto_625(I_2821_D, I_2855_S);
	nand auto_626(I_2853_S, I_2791_S, I_3241_D);
	nor auto_627(I_2794_D, I_3271_S, I_2951_S, I_3111_S);
	not auto_628(I_2735_D, I_3019_S);
	not auto_629(I_2741_D, I_2869_D);
	not auto_630(I_2745_D, I_2713_D);
	not auto_631(I_2747_D, I_1755_D);
	not auto_632(I_2749_D, I_2009_D);
	nand auto_633(I_2815_D, I_2559_S, I_2718_S, I_2157_S);
	nand auto_634(I_2855_S, I_2853_D, I_3241_D);
	nand auto_635(I_277_D, I_341_D, I_341_D);
	not auto_636(I_2775_D, I_2711_S);
	not auto_637(I_2809_D, I_2745_D); // NMOS strength = 2
	nand auto_638(I_2811_D, I_1755_D, I_2649_D);
	nand auto_639(I_2813_D, I_2875_D, I_2009_D);
	not auto_640(I_2817_D, I_2753_D);
	not auto_641(I_2791_S, I_2855_D);
	not auto_642(I_2799_S, I_3823_S);
	not auto_643(I_2805_S, I_2709_S);
	not auto_644(I_2807_S, I_2775_D);
	nand auto_645(I_2955_D, I_3751_S, I_3271_S, I_2951_S, I_3111_S);
	not auto_646(I_315_D, I_251_S); // NMOS strength = 2
	nand auto_647(I_2865_D, I_1679_D, I_3116_D);
	nand auto_648(I_2875_D, I_2811_D, I_2715_D);
	nand auto_649(I_2877_D, I_2749_D, I_3133_D);
	not auto_650(I_2879_D, I_2717_D); // NMOS strength = 2
	nand auto_651(I_3169_S, I_2881_G, I_2945_S);
	not auto_652(I_2981_D, I_3015_S);
	nand auto_653(I_3013_S, I_3241_D, I_2951_S);
	not auto_654(I_2889_D, I_1033_D);
	not auto_655(I_2893_D, I_2253_D);
	nor auto_656(I_2928_D, I_1679_D, I_3116_D);
	not auto_657(I_93_S, I_503_G); // NMOS strength = 3
	not auto_658(I_2905_D, I_2873_D);
	not auto_659(I_2907_D, I_1755_D);
	nand auto_660(I_2972_D, I_2877_D, I_2813_D);
	nand auto_661(I_2975_D, I_3198_S, I_3036_G, I_3038_S);
	nand auto_662(I_3015_S, I_3241_D, I_3013_D);
	nand auto_663(I_2953_D, I_2955_D, I_1033_D);
	nand auto_664(I_2957_D, I_3339_D, I_2253_D);
	not auto_665(I_2969_D, I_2905_D); // NMOS strength = 2
	nand auto_666(I_2971_D, I_2809_D, I_1755_D);
	not auto_667(I_2945_S, I_3009_D);
	not auto_668(I_2951_S, I_3015_D);
	not auto_669(I_2961_S, I_2928_D);
	not auto_670(I_297_S, I_616_S);
	nand auto_671(I_3075_D, I_2632_D, I_2791_S, I_3173_S, I_3171_D);
	nand auto_672(I_3017_D, I_2889_D, I_3083_D);
	nand auto_673(I_3021_D, I_3271_S, I_2893_D);
	nand auto_674(I_3023_D, I_3116_D, I_3019_S);
	not auto_675(I_3_D, I_3_G);
	nand auto_676(I_3035_D, I_3031_D, I_2907_D);
	not auto_677(I_3036_S, I_3036_G);
	not auto_678(I_3038_S, I_1597_D);
	not auto_679(I_3019_S, I_3019_G);
	not auto_680(I_3039_S, I_3038_S);
	nand auto_681(I_3073_D, I_3073_G, I_3169_D);
	not auto_682(I_3141_D, I_3175_S);
	nand auto_683(I_3173_S, I_3111_S, I_3241_D);
	nand auto_684(I_3112_D, I_2953_D, I_3017_D);
	nand auto_685(I_3083_D, I_3657_D, I_2951_S);
	nand auto_686(I_3116_D, I_2957_D, I_3021_D);
	nor auto_687(I_3086_D, I_3116_D, I_3019_S);
	nand auto_688(I_3345_S, I_2961_S, I_2865_D);
	not auto_689(I_3059_D, I_3219_D);
	not auto_690(I_3061_D, I_3191_S);
	not auto_691(I_3063_D, I_3191_D);
	not auto_692(I_3065_D, I_3033_D);
	nand auto_693(I_3130_D, I_3035_D, I_2971_D);
	nand auto_694(I_3133_D, I_3135_D, I_2975_D, I_3295_D);
	nand auto_695(I_3135_D, I_3659_S, I_3038_S, I_3199_S);
	nand auto_696(I_3175_S, I_3241_D, I_3173_D);
	not auto_697(I_3129_D, I_3065_D); // NMOS strength = 2
	not auto_698(I_95_D, I_95_G); // NMOS strength = 3
	not auto_699(I_3137_D, I_3073_D);
	not auto_700(I_3111_S, I_3175_D);
	not auto_701(I_3119_S, I_3086_D);
	not auto_702(I_3313_D, I_3345_S);
	not auto_703(I_3123_S, I_3985_D);
	not auto_704(I_3125_S, I_3345_D);
	not auto_705(I_3127_S, I_3031_S);
	nand auto_706(I_3171_D, I_3173_S, I_3013_S);
	nand auto_707(I_3177_D, I_1283_D, I_3112_D);
	nand auto_708(I_3193_D, I_3449_D, I_3225_D);
	nand auto_709(I_3197_D, I_3453_D, I_3229_D);
	not auto_710(I_3198_S, I_1821_D);
	not auto_711(I_3195_S, I_3195_G);
	not auto_712(I_3199_S, I_3198_S);
	nand auto_713(I_3489_S, I_3201_G, I_3265_S);
	not auto_714(I_3301_D, I_3335_S);
	nand auto_715(I_3333_S, I_3271_S, I_3241_D);
	not auto_716(I_3241_D, I_3177_D); // NMOS strength = 2
	not auto_717(I_321_D, I_33_D);
	nand auto_718(I_3503_S, I_3119_S, I_3023_D);
	nand auto_719(I_3287_D, I_3510_S, I_3347_D, I_3350_S);
	not auto_720(I_3225_D, I_1689_D);
	nand auto_721(I_3291_D, VDD, I_3514_S, I_3354_S);
	not auto_722(I_3229_D, I_2009_D);
	nand auto_723(I_355_D, I_1029_D, I_1249_D);
	nand auto_724(I_3295_D, I_3039_S, I_3198_S, VSS);
	nand auto_725(I_3335_S, I_3333_D, I_3241_D);
	not auto_726(I_3249_D, I_3185_S);
	nand auto_727(I_421_D, I_1187_S, I_389_S);
	nand auto_728(I_3285_D, I_3413_D, I_3349_D);
	nand auto_729(I_3289_D, I_1689_D, I_3285_D);
	nand auto_730(I_3293_D, I_2009_D, I_3130_D);
	not auto_731(I_3265_S, I_3329_D);
	not auto_732(I_423_D, I_453_S);
	not auto_733(I_3271_S, I_3335_D);
	not auto_734(I_3471_D, I_3503_S);
	not auto_735(I_3281_S, I_3249_D);
	not auto_736(I_3283_S, I_3189_S);
	not auto_737(I_329_D, I_395_D);
	not auto_738(I_3331_D, I_3331_G); // NMOS strength = 2
	nand auto_739(I_395_D, I_297_S, I_618_S, I_461_S);
	nand auto_740(I_3349_D, I_1831_S, I_3445_S);
	not auto_741(I_3350_S, I_1597_D);
	nand auto_742(I_3353_D, I_3193_D, I_3289_D);
	not auto_743(I_3354_S, I_1597_D);
	nand auto_744(I_3357_D, I_3293_D, I_3197_D);
	not auto_745(I_3359_D, I_2972_D); // NMOS strength = 2
	not auto_746(I_3351_S, I_3350_S);
	not auto_747(I_3355_S, I_3354_S);
	nand auto_748(I_3393_D, I_3489_D, I_3393_G);
	not auto_749(I_3363_D, I_3491_S);
	not auto_750(I_3461_D, I_3495_S);
	nand auto_751(I_3493_S, I_3431_S, I_3241_D);
	not auto_752(I_3369_D, I_3591_S);
	not auto_753(I_3371_D, I_3499_D);
	not auto_754(I_3379_D, I_3507_D);
	nand auto_755(I_3413_D, I_3381_G, I_3735_G);
	nand auto_756(I_3447_D, I_3987_S, I_3350_S, I_3511_S);
	nand auto_757(I_3449_D, I_3447_D, I_3287_D, I_3607_D);
	nand auto_758(I_3451_D, I_3354_S, I_3983_D, I_3515_S);
	nand auto_759(I_3453_D, I_3291_D, I_3451_D, I_3611_D);
	not auto_760(I_3423_D, I_3357_D); // NMOS strength = 2
	nand auto_761(I_3427_D, I_2853_S, I_3013_S);
	nand auto_762(I_3495_S, I_3241_D, I_3493_D);
	nand auto_763(I_3663_S, I_3501_D, I_3565_D);
	not auto_764(I_3407_D, I_3535_D);
	nand auto_765(I_341_D, I_437_D, I_437_D);
	not auto_766(I_3457_D, I_3393_D);
	not auto_767(I_375_D, I_471_D); // NMOS strength = 2
	not auto_768(I_3431_S, I_3495_D);
	not auto_769(I_3433_S, I_3499_D);
	not auto_770(I_3435_S, I_3497_S);
	not auto_771(I_3439_S, I_3407_D);
	not auto_772(I_3443_S, I_3503_D);
	not auto_773(I_3445_S, I_3735_G);
	not auto_774(I_443_D, I_313_D); // NMOS strength = 2
	nand auto_775(I_3501_D, I_3431_S, I_3597_S);
	not auto_776(I_347_D, I_603_D);
	nand auto_777(I_3505_D, I_2319_D, I_3663_S);
	not auto_778(I_3510_S, I_1821_D);
	not auto_779(I_3514_S, I_1821_D);
	nand auto_780(I_3517_D, I_3773_D, I_3549_D);
	not auto_781(I_3519_D, I_3677_D); // NMOS strength = 2
	not auto_782(I_477_S, I_317_D);
	nor auto_783(I_3491_S, I_3587_D, I_3427_D);
	nand auto_784(I_447_D, I_639_S, I_319_D);
	not auto_785(I_3511_S, I_3510_S);
	not auto_786(I_3515_S, I_3514_S);
	not auto_787(I_3521_D, I_3555_G);
	nand auto_788(I_3587_D, I_3555_G, I_3333_S, I_3173_S);
	not auto_789(I_3621_D, I_3655_S);
	nand auto_790(I_3653_S, I_3241_D, I_3591_S);
	not auto_791(I_3529_D, I_3529_G);
	not auto_792(I_385_D, I_448_D); // NMOS strength = 2
	nor auto_793(I_3562_D, I_3657_D, I_3431_S);
	nand auto_794(I_3565_D, I_2253_D, I_3499_S);
	not auto_795(I_3535_D, I_3599_S);
	nor auto_796(I_3568_D, I_3663_S, I_2319_D);
	nand auto_797(I_3607_D, I_3351_S, I_3510_S, I_1962_D);
	nand auto_798(I_3609_D, I_3027_D, I_3832_S, I_3672_S);
	nand auto_799(I_3611_D, I_3355_S, I_3514_S, VDD);
	not auto_800(I_3549_D, I_1689_D);
	nand auto_801(I_3615_D, I_3029_D, I_3838_S, I_3678_S);
	nand auto_802(I_3585_D, I_3975_D, I_3913_S);
	nand auto_803(I_3655_S, I_3241_D, I_3653_D);
	nand auto_804(I_3613_D, I_1689_D, I_3997_D);
	nand auto_805(I_453_S, I_1187_S, I_455_D);
	not auto_806(I_3593_S, I_3593_G);
	not auto_807(I_3595_S, I_3593_S);
	not auto_808(I_3597_S, I_2253_D);
	not auto_809(I_3599_S, I_3825_D);
	not auto_810(I_3601_S, I_3568_D);
	not auto_811(I_3649_D, I_3649_G); // NMOS strength = 2
	not auto_812(I_3651_D, I_3755_S); // NMOS strength = 2
	not auto_813(I_3657_D, I_3813_S); // NMOS strength = 2
	nand auto_814(I_3725_D, I_3595_S, I_3919_S, I_3691_D, I_3859_D);
	not auto_815(I_3672_S, I_1597_D);
	not auto_816(I_3675_D, I_3995_D); // NMOS strength = 2
	nand auto_817(I_3677_D, I_3517_D, I_3613_D);
	not auto_818(I_3678_S, I_1597_D);
	not auto_819(I_3659_S, I_3659_G);
	not auto_820(I_3673_S, I_3672_S);
	not auto_821(I_3679_S, I_3678_S);
	not auto_822(I_3681_D, I_3649_D);
	not auto_823(I_3683_D, I_3649_D);
	not auto_824(I_3781_D, I_3815_S);
	nand auto_825(I_3813_S, I_3241_D, I_3751_S);
	nand auto_826(I_3753_D, I_3969_S, I_3915_G, I_3847_G);
	not auto_827(I_3691_D, I_3659_S);
	not auto_828(I_3695_D, I_3823_D);
	nand auto_829(I_3985_S, I_3601_S, I_3505_D);
	not auto_830(I_3699_D, I_3827_D);
	nand auto_831(I_101_D, I_69_S, I_1187_S);
	not auto_832(I_3701_D, I_3829_D);
	not auto_833(I_3703_D, I_3735_G);
	nand auto_834(I_3769_D, I_3990_S, I_3672_S, I_3833_S);
	nand auto_835(I_3771_D, I_3609_D, I_3769_D, I_3929_D);
	nand auto_836(I_3773_D, I_3775_D, I_3615_D, I_3935_D);
	nand auto_837(I_3775_D, I_3988_S, I_3678_S, I_3839_S);
	nand auto_838(I_3745_D, I_3649_D, I_2791_S);
	nand auto_839(I_3747_D, I_1741_S, I_3649_D);
	nand auto_840(I_3815_S, I_3241_D, I_3813_D);
	nand auto_841(I_3767_D, I_3767_G, I_3735_G);
	not auto_842(I_3751_S, I_3815_D);
	nor auto_843(I_3755_S, I_3883_D, I_3725_D);
	not auto_844(I_3759_S, I_3663_S);
	not auto_845(I_3953_D, I_3985_S);
	not auto_846(I_3763_S, I_3667_S);
	not auto_847(I_3765_S, I_3669_S);
	nand auto_848(I_3809_D, I_3681_D, I_2631_S);
	nand auto_849(I_3811_D, I_3683_D, I_2791_S);
	nand auto_850(I_3817_D, I_3847_D, I_3977_G);
	nand auto_851(I_3883_D, I_3988_S, I_3819_G, I_3851_G, I_3887_D);
	nand auto_852(I_3831_D, I_3830_G, I_3703_D);
	not auto_853(I_3832_S, I_1821_D);
	nand auto_854(I_3835_D, I_3867_D, I_3771_D);
	nand auto_855(I_3837_D, I_3869_D, I_3836_G);
	not auto_856(I_3838_S, I_1821_D);
	not auto_857(I_3833_S, I_3832_S);
	not auto_858(I_3839_S, I_3838_S);
	nand auto_859(I_3904_D, I_3745_D, I_3809_D);
	nand auto_860(I_3906_D, I_3747_D, I_3811_D);
	not auto_861(I_3845_D, I_3649_D);
	not auto_862(I_3847_D, I_3847_G);
	nand auto_863(I_3913_S, I_3753_D, I_3817_D, I_3977_D);
	not auto_864(I_3859_D, I_3923_S);
	not auto_865(I_3861_D, I_3195_S);
	nand auto_866(I_3926_D, I_3767_D, I_3831_D);
	nand auto_867(I_3929_D, I_3673_S, I_3832_S, I_3129_D);
	not auto_868(I_3867_D, I_1689_D);
	not auto_869(I_3869_D, I_1755_D);
	not auto_870(I_387_S, I_1249_D);
	nand auto_871(I_3935_D, I_3679_S, I_3838_S, I_2969_D);
	nand auto_872(I_3909_D, I_3649_D, I_2631_S);
	nand auto_873(I_3911_D, I_3845_D, I_3911_G);
	not auto_874(I_3887_D, I_3987_S);
	not auto_875(I_3889_D, I_3825_S);
	not auto_876(I_389_S, I_453_D);
	nand auto_877(I_3931_D, I_1689_D, I_3926_D);
	nand auto_878(I_133_S, I_1187_S, I_135_D);
	nand auto_879(I_3933_D, I_1755_D, I_3933_G);
	not auto_880(I_3915_S, I_3915_G);
	not auto_881(I_3917_S, I_3529_D);
	not auto_882(I_3919_S, I_3983_D);
	not auto_883(I_3921_S, I_3889_D);
	not auto_884(I_3923_S, I_3923_G);
	not auto_885(I_393_S, I_555_D);
	nand auto_886(I_3973_D, I_3911_D, I_3909_D);
	nand auto_887(I_3975_D, I_3755_S, I_3974_G);
	nand auto_888(I_3977_D, I_3977_G, I_3915_S);
	not auto_889(I_3979_D, I_3981_D); // NMOS strength = 2
	nand auto_890(I_3981_D, I_3917_S, I_3980_G);
	not auto_891(I_3983_D, I_3982_G);
	not auto_892(I_3988_S, I_3988_G);
	not auto_893(I_3990_S, I_3990_G);
	nand auto_894(I_3995_D, I_3931_D, I_3835_D);
	nand auto_895(I_3997_D, I_3933_D, I_3837_D);
	not auto_896(I_3999_D, I_3999_G); // NMOS strength = 2
	not auto_897(I_3969_S, I_3971_S);
	not auto_898(I_3971_S, I_3971_G);
	not auto_899(I_3987_S, I_3987_G);
	not auto_900(I_3993_S, I_3993_G);
	not auto_901(I_439_D, I_375_D);
	not auto_902(I_409_S, I_443_D);
	not auto_903(I_445_D, I_477_S);
	not auto_904(I_415_S, I_447_D);
	nor auto_905(I_448_D, I_1089_D, I_545_D);
	nand auto_906(I_457_D, I_3065_D, I_2905_D);
	not auto_907(I_458_S, I_461_S);
	nand auto_908(I_437_D, I_1373_S, I_1373_S);
	not auto_909(I_461_S, I_2809_D);
	nand auto_910(I_581_D, I_549_S, I_1187_S);
	not auto_911(I_583_D, I_613_S);
	nand auto_912(I_553_D, I_524_D, I_3065_D, I_2905_D);
	nand auto_913(I_555_D, I_458_S, I_616_S, I_618_S);
	nor auto_914(I_524_D, I_493_G, I_1211_D);
	not auto_915(I_503_D, I_503_G);
	not auto_916(I_505_D, I_601_D);
	not auto_917(I_2201_D, I_507_G);
	not auto_918(I_509_D, I_573_D);
	not auto_919(I_511_D, I_479_D);
	nand auto_920(I_545_D, I_609_D, auto_net_3);
	or auto_921(auto_net_3, I_1832_D, I_547_D);
	nand auto_922(I_547_D, I_611_D, I_675_D);
	nand auto_923(I_613_S, I_1187_S, I_615_D);
	not auto_924(I_601_D, I_473_D); // NMOS strength = 2
	nand auto_925(I_573_D, I_511_D, I_957_S);
	not auto_926(I_549_S, I_613_D);
	not auto_927(I_2841_D, I_571_G);
	not auto_928(I_575_S, I_511_D);
	nand auto_929(I_609_D, I_1832_D, I_547_D);
	nand auto_930(I_611_D, I_707_S, I_709_S);
	not auto_931(I_616_S, I_2649_D);
	not auto_932(I_618_S, I_553_D);
	nand auto_933(I_603_D, I_667_D, I_667_D);
	nand auto_934(I_675_D, I_1189_D, I_1249_D);
	nand auto_935(I_741_D, I_1187_S, I_709_S);
	not auto_936(I_743_D, I_773_S);
	not auto_937(I_65_S, I_128_D);
	nand auto_938(I_715_D, I_616_S, I_461_S, I_618_S);
	not auto_939(I_759_D, I_727_D);
	not auto_940(I_763_D, I_633_D); // NMOS strength = 2
	nand auto_941(I_667_D, I_827_D, I_827_D);
	nand auto_942(I_765_D, I_637_D, I_799_S);
	nor auto_943(I_67_S, I_3_D, I_65_S);
	not auto_944(I_705_D, I_768_D); // NMOS strength = 2
	nand auto_945(I_773_S, I_1187_S, I_775_D);
	not auto_946(I_69_S, I_133_D);
	not auto_947(I_727_D, I_791_D); // NMOS strength = 2
	not auto_948(I_103_D, I_133_S);
	not auto_949(I_735_D, I_575_S); // NMOS strength = 2
	not auto_950(I_707_S, I_1249_D);
	not auto_951(I_709_S, I_773_D);
	not auto_952(I_713_S, I_235_D);
	not auto_953(I_789_D, I_1045_D); // NMOS strength = 3
	not auto_954(I_729_S, I_763_D);
	not auto_955(I_733_S, I_765_D);
	nor auto_956(I_768_D, I_1089_D, I_865_D);
	not auto_957(I_779_S, I_713_S);
	nand auto_958(I_901_D, I_869_S, I_1187_S);
	not auto_959(I_903_D, I_933_S);
	not auto_960(I_809_D, I_777_D);
	nand auto_961(I_821_D, I_917_D, I_917_D);
	not auto_962(I_855_D, I_951_D); // NMOS strength = 2
	not auto_963(I_825_D, I_921_D);
	nand auto_964(I_827_D, I_923_D, I_923_D);
	not auto_965(I_957_S, I_797_D);
	nand auto_966(I_1439_S, I_415_S, I_733_S, I_1055_S);
	nand auto_967(I_865_D, I_929_D, auto_net_4);
	or auto_968(auto_net_4, I_1832_D, I_867_D);
	nand auto_969(I_867_D, I_995_D, I_931_D);
	nand auto_970(I_933_S, I_935_D, I_1187_S);
	not auto_971(I_873_D, I_809_D); // NMOS strength = 2
	not auto_972(I_2681_D, I_85_G);
	not auto_973(I_921_D, I_793_D); // NMOS strength = 2
	not auto_974(I_869_S, I_933_D);
	not auto_975(I_2361_D, I_87_G);
	not auto_976(I_919_D, I_855_D);
	not auto_977(I_925_D, I_957_S);
	nand auto_978(I_929_D, I_867_D, I_1832_D);
	nand auto_979(I_931_D, I_1027_S, I_869_S);
	not auto_980(I_2041_D, I_91_G);
	nand auto_981(I_917_D, I_1331_D, I_1331_D);
	nand auto_982(I_923_D, I_989_D, I_989_D);
	nand auto_983(I_995_D, I_1349_D, I_1249_D);
	not auto_984(I_1061_D, I_1029_D);
	nand auto_985(I_1063_D, I_1093_S, I_1187_S);
	not auto_986(I_969_D, I_937_D);
	nor auto_987(I_128_D, I_1089_D, I_225_D);
	not auto_988(I_975_D, I_1997_D);
	nand auto_989(I_983_D, I_1113_S, I_1113_S);
	not auto_990(I_989_D, I_511_D);
	generic_pmos I_1393(.D(I_1393_D), .G(I_1361_S), .S(I_1999_D));
	generic_nmos I_1424(.D(I_1425_S), .G(I_1361_S), .S(VSS));
	generic_nmos I_1654(.D(VSS), .G(I_151_D), .S(VSS));
	generic_pmos I_1655(.D(VDD), .G(I_151_D), .S(VDD));
	generic_nmos I_1712(.D(VSS), .G(I_1648_D), .S(I_2545_S));
	generic_nmos I_1714(.D(VSS), .G(I_2133_G), .S(VSS));
	generic_pmos I_1745(.D(I_2545_S), .G(I_1585_D), .S(VDD));
	generic_pmos I_1747(.D(VDD), .G(I_2133_G), .S(VDD));
	generic_nmos I_1966(.D(VSS), .G(I_2063_D), .S(I_1998_D));
	generic_pmos I_1967(.D(VDD), .G(I_2063_D), .S(I_1999_D));
	generic_nmos I_1998(.D(I_1998_D), .G(I_2127_D), .S(I_1999_D));
	generic_pmos I_1999(.D(I_1999_D), .G(I_2127_D), .S(VDD));
	generic_nmos I_2196(.D(VSS), .G(I_2132_D), .S(I_2711_S));
	generic_pmos I_2199(.D(I_2199_D), .G(I_2167_S), .S(I_2231_D));
	generic_pmos I_2229(.D(I_2711_S), .G(I_2069_D), .S(VDD));
	generic_nmos I_2230(.D(I_2231_S), .G(I_2167_S), .S(VSS));
	generic_nmos I_2250(.D(I_3499_D), .G(I_873_D), .S(I_2282_D));
	generic_pmos I_2251(.D(VDD), .G(I_873_D), .S(I_3499_D));
	generic_nmos I_2282(.D(I_2282_D), .G(I_2219_S), .S(VSS));
	generic_pmos I_2283(.D(I_3499_D), .G(I_2219_S), .S(VDD));
	generic_pmos I_2349(.D(VDD), .G(I_3337_D), .S(VDD));
	generic_nmos I_2352(.D(VSS), .G(I_2288_D), .S(I_3185_S));
	generic_nmos I_2380(.D(VSS), .G(I_3337_D), .S(VSS));
	generic_pmos I_2385(.D(I_3185_S), .G(I_2225_D), .S(VDD));
	generic_nmos I_2508(.D(VSS), .G(I_3591_S), .S(VSS));
	generic_nmos I_2518(.D(VSS), .G(I_2454_D), .S(I_2869_D));
	generic_pmos I_2541(.D(VDD), .G(I_3591_S), .S(VDD));
	generic_pmos I_2551(.D(I_2869_D), .G(I_2391_D), .S(VDD));
	generic_nmos I_2768(.D(VSS), .G(I_3065_D), .S(VSS));
	generic_pmos I_2769(.D(VDD), .G(I_3065_D), .S(VDD));
	generic_nmos I_2802(.D(VSS), .G(I_2709_S), .S(VSS));
	generic_pmos I_2803(.D(VDD), .G(I_2709_S), .S(VDD));
	generic_pmos I_2837(.D(I_2837_D), .G(I_2805_S), .S(I_2869_D));
	generic_nmos I_2868(.D(I_3191_D), .G(I_2805_S), .S(VSS));
	generic_nmos I_2992(.D(VSS), .G(I_2928_D), .S(I_3825_S));
	generic_pmos I_3025(.D(I_3825_S), .G(I_2865_D), .S(VDD));
	generic_pmos I_3149(.D(I_3149_D), .G(I_3593_S), .S(I_3181_D));
	generic_nmos I_3150(.D(VSS), .G(I_3086_D), .S(I_3823_D));
	generic_pmos I_3155(.D(I_3155_D), .G(I_3123_S), .S(I_3219_D));
	generic_pmos I_3157(.D(I_3157_D), .G(I_3125_S), .S(I_3191_S));
	generic_pmos I_3159(.D(I_3159_D), .G(I_3127_S), .S(I_3191_D));
	generic_nmos I_3180(.D(I_3180_D), .G(I_3593_S), .S(I_3180_S));
	generic_pmos I_3183(.D(I_3823_D), .G(I_3023_D), .S(VDD));
	generic_nmos I_3186(.D(I_3507_D), .G(I_3123_S), .S(VSS));
	generic_nmos I_3188(.D(I_3189_S), .G(I_3125_S), .S(VSS));
	generic_nmos I_3190(.D(I_3191_S), .G(I_3127_S), .S(VSS));
	generic_nmos I_3218(.D(I_3219_D), .G(I_3283_S), .S(VSS));
	generic_pmos I_3219(.D(I_3219_D), .G(I_3283_S), .S(VDD));
	generic_nmos I_3372(.D(VSS), .G(I_3659_S), .S(VSS));
	generic_pmos I_3373(.D(VDD), .G(I_3659_S), .S(VDD));
	generic_pmos I_3465(.D(I_3465_D), .G(I_3433_S), .S(I_3591_S));
	generic_pmos I_3467(.D(I_3467_D), .G(I_3435_S), .S(I_3499_D));
	generic_pmos I_3475(.D(I_3475_D), .G(I_3443_S), .S(I_3507_D));
	generic_nmos I_3496(.D(I_3497_S), .G(I_3433_S), .S(VSS));
	generic_nmos I_3498(.D(I_3499_S), .G(I_3435_S), .S(VSS));
	generic_nmos I_3506(.D(I_3827_D), .G(I_3443_S), .S(VSS));
	generic_nmos I_3590(.D(VSS), .G(I_3655_D), .S(I_3591_S));
	generic_pmos I_3591(.D(VDD), .G(I_3655_D), .S(I_3591_S));
	generic_nmos I_3632(.D(VSS), .G(I_3568_D), .S(I_3825_D));
	generic_pmos I_3665(.D(I_3825_D), .G(I_3505_D), .S(VDD));
	generic_nmos I_3756(.D(VSS), .G(I_3659_S), .S(I_3788_D));
	generic_pmos I_3757(.D(VDD), .G(I_3659_S), .S(I_3884_D));
	generic_nmos I_3788(.D(I_3788_D), .G(I_3983_D), .S(I_3820_D));
	generic_pmos I_3789(.D(VDD), .G(I_3977_G), .S(I_3884_D));
	generic_pmos I_3791(.D(I_3791_D), .G(I_3759_S), .S(I_3823_D));
	generic_pmos I_3795(.D(I_3795_D), .G(I_3763_S), .S(I_3827_D));
	generic_pmos I_3797(.D(I_3797_D), .G(I_3765_S), .S(I_3829_D));
	generic_nmos I_3820(.D(I_3820_D), .G(I_3977_G), .S(I_3852_D));
	generic_pmos I_3821(.D(I_3884_D), .G(I_3983_D), .S(VDD));
	generic_nmos I_3822(.D(I_3823_S), .G(I_3759_S), .S(VSS));
	generic_nmos I_3826(.D(I_3829_D), .G(I_3763_S), .S(VSS));
	generic_nmos I_3828(.D(I_3829_S), .G(I_3765_S), .S(VSS));
	generic_nmos I_3852(.D(I_3852_D), .G(I_3529_D), .S(I_3884_D));
	generic_pmos I_3853(.D(I_3884_D), .G(I_3529_D), .S(VDD));
	generic_nmos I_3884(.D(I_3884_D), .G(VSS), .S(VSS));
	generic_pmos I_3885(.D(VDD), .G(VSS), .S(VDD));
	generic_nmos I_3890(.D(VSS), .G(I_3861_D), .S(VSS));
	generic_pmos I_3891(.D(VDD), .G(I_3861_D), .S(VDD));
	generic_cmos pass_1(.gn(I_329_D), .gp(I_395_D), .p1(I_101_D), .p2(I_133_D));
	generic_cmos pass_10(.gn(I_93_S), .gp(I_95_D), .p1(I_1117_D), .p2(I_1407_D));
	generic_cmos pass_100(.gn(I_2053_S), .gp(I_1991_S), .p1(I_2181_D), .p2(I_2213_D));
	generic_cmos pass_101(.gn(I_1991_S), .gp(I_2053_S), .p1(I_2213_S), .p2(I_2215_D));
	generic_cmos pass_102(.gn(I_1973_D), .gp(I_2007_D), .p1(I_2201_D), .p2(I_2233_D));
	generic_cmos pass_103(.gn(I_2305_S), .gp(I_2529_S), .p1(I_2209_D), .p2(I_2209_S));
	generic_cmos pass_104(.gn(I_1991_S), .gp(I_2053_S), .p1(I_2213_D), .p2(I_2213_S));
	generic_cmos pass_105(.gn(I_2053_S), .gp(I_1991_S), .p1(I_2215_D), .p2(I_2215_S));
	generic_cmos pass_106(.gn(I_2071_S), .gp(I_2167_S), .p1(I_2231_D), .p2(I_2231_S));
	generic_cmos pass_107(.gn(I_2007_D), .gp(I_1973_D), .p1(I_2233_D), .p2(I_2329_D));
	generic_cmos pass_108(.gn(I_2625_S), .gp(I_2657_D), .p1(I_2529_S), .p2(I_2369_D));
	generic_cmos pass_109(.gn(I_2213_S), .gp(I_2151_S), .p1(I_2341_D), .p2(I_2373_D));
	generic_cmos pass_11(.gn(I_93_S), .gp(I_95_D), .p1(I_1119_D), .p2(I_1247_D));
	generic_cmos pass_110(.gn(I_2151_S), .gp(I_2213_S), .p1(I_2373_S), .p2(I_2375_D));
	generic_cmos pass_111(.gn(I_1973_D), .gp(I_2007_D), .p1(I_2361_D), .p2(I_2393_D));
	generic_cmos pass_112(.gn(I_2657_D), .gp(I_2625_S), .p1(I_2369_D), .p2(I_2433_D));
	generic_cmos pass_113(.gn(I_2151_S), .gp(I_2213_S), .p1(I_2373_D), .p2(I_2373_S));
	generic_cmos pass_114(.gn(I_2213_S), .gp(I_2151_S), .p1(I_2375_D), .p2(I_2375_S));
	generic_cmos pass_115(.gn(I_2517_D), .gp(I_2549_S), .p1(I_2711_S), .p2(I_2389_S));
	generic_cmos pass_116(.gn(I_2007_D), .gp(I_1973_D), .p1(I_2393_D), .p2(I_2489_D));
	generic_cmos pass_117(.gn(I_2657_D), .gp(I_2625_S), .p1(I_2497_D), .p2(I_2529_D));
	generic_cmos pass_118(.gn(I_2530_S), .gp(I_2535_G), .p1(I_2501_D), .p2(I_2533_D));
	generic_cmos pass_119(.gn(I_2535_G), .gp(I_2534_G), .p1(I_2533_S), .p2(I_2535_D));
	generic_cmos pass_12(.gn(I_315_D), .gp(I_251_S), .p1(I_155_D), .p2(I_153_D));
	generic_cmos pass_120(.gn(I_2453_D), .gp(I_2485_S), .p1(I_2517_D), .p2(I_2549_D));
	generic_cmos pass_121(.gn(I_1973_D), .gp(I_2007_D), .p1(I_2521_D), .p2(I_2553_D));
	generic_cmos pass_122(.gn(I_2625_S), .gp(I_2657_D), .p1(I_2529_D), .p2(I_2529_S));
	generic_cmos pass_123(.gn(I_2535_G), .gp(I_2534_G), .p1(I_2533_D), .p2(I_2533_S));
	generic_cmos pass_124(.gn(I_2534_G), .gp(I_2535_G), .p1(I_2535_D), .p2(I_2535_S));
	generic_cmos pass_125(.gn(I_2673_D), .gp(I_2705_S), .p1(I_3185_S), .p2(I_2545_S));
	generic_cmos pass_126(.gn(I_2485_S), .gp(I_2453_D), .p1(I_2549_D), .p2(I_2549_S));
	generic_cmos pass_127(.gn(I_2007_D), .gp(I_1973_D), .p1(I_2553_D), .p2(I_2649_D));
	generic_cmos pass_128(.gn(I_329_D), .gp(I_395_D), .p1(I_261_D), .p2(I_293_D));
	generic_cmos pass_129(.gn(I_395_D), .gp(I_329_D), .p1(I_263_D), .p2(I_295_D));
	generic_cmos pass_13(.gn(I_1097_S), .gp(I_715_D), .p1(I_1221_D), .p2(I_1253_D));
	generic_cmos pass_130(.gn(I_2945_S), .gp(I_3169_S), .p1(I_2657_D), .p2(I_2689_D));
	generic_cmos pass_131(.gn(I_2533_S), .gp(I_2471_S), .p1(I_2661_D), .p2(I_2693_D));
	generic_cmos pass_132(.gn(I_2471_S), .gp(I_2533_S), .p1(I_2693_S), .p2(I_2695_D));
	generic_cmos pass_133(.gn(I_2799_S), .gp(I_3823_S), .p1(I_3019_S), .p2(I_3669_S));
	generic_cmos pass_134(.gn(I_2609_D), .gp(I_2641_S), .p1(I_2673_D), .p2(I_3031_S));
	generic_cmos pass_135(.gn(I_2869_D), .gp(I_2741_D), .p1(I_2805_S), .p2(I_2709_D));
	generic_cmos pass_136(.gn(I_1973_D), .gp(I_2007_D), .p1(I_2681_D), .p2(I_2713_D));
	generic_cmos pass_137(.gn(I_3169_S), .gp(I_2945_S), .p1(I_2689_D), .p2(I_2753_D));
	generic_cmos pass_138(.gn(I_2471_S), .gp(I_2533_S), .p1(I_2693_D), .p2(I_2693_S));
	generic_cmos pass_139(.gn(I_2533_S), .gp(I_2471_S), .p1(I_2695_D), .p2(I_2695_S));
	generic_cmos pass_14(.gn(I_715_D), .gp(I_1097_S), .p1(I_1223_D), .p2(I_1255_D));
	generic_cmos pass_140(.gn(I_3823_S), .gp(I_2799_S), .p1(I_3669_S), .p2(I_2735_D));
	generic_cmos pass_141(.gn(I_2641_S), .gp(I_2609_D), .p1(I_3031_S), .p2(I_2705_S));
	generic_cmos pass_142(.gn(I_2741_D), .gp(I_2869_D), .p1(I_2709_D), .p2(I_2709_S));
	generic_cmos pass_143(.gn(I_2839_D), .gp(I_2871_S), .p1(I_2869_D), .p2(I_2711_S));
	generic_cmos pass_144(.gn(I_2007_D), .gp(I_1973_D), .p1(I_2713_D), .p2(I_2809_D));
	generic_cmos pass_145(.gn(I_315_D), .gp(I_251_S), .p1(I_279_D), .p2(I_311_D));
	generic_cmos pass_146(.gn(I_251_S), .gp(I_315_D), .p1(I_281_D), .p2(I_313_D));
	generic_cmos pass_147(.gn(I_3169_S), .gp(I_2945_S), .p1(I_2817_D), .p2(I_2849_D));
	generic_cmos pass_148(.gn(I_2693_S), .gp(I_2631_S), .p1(I_2821_D), .p2(I_2853_D));
	generic_cmos pass_149(.gn(I_2631_S), .gp(I_2693_S), .p1(I_2853_S), .p2(I_2855_D));
	generic_cmos pass_15(.gn(I_1258_G), .gp(I_1099_S), .p1(I_1225_D), .p2(I_1257_D));
	generic_cmos pass_150(.gn(I_2775_D), .gp(I_2807_S), .p1(I_2839_D), .p2(I_2871_D));
	generic_cmos pass_151(.gn(I_1973_D), .gp(I_2007_D), .p1(I_2841_D), .p2(I_2873_D));
	generic_cmos pass_152(.gn(I_2945_S), .gp(I_3169_S), .p1(I_2849_D), .p2(I_2849_S));
	generic_cmos pass_153(.gn(I_95_D), .gp(I_93_S), .p1(I_285_D), .p2(I_317_D));
	generic_cmos pass_154(.gn(I_2631_S), .gp(I_2693_S), .p1(I_2853_D), .p2(I_2853_S));
	generic_cmos pass_155(.gn(I_2693_S), .gp(I_2631_S), .p1(I_2855_D), .p2(I_2855_S));
	generic_cmos pass_156(.gn(I_2709_S), .gp(I_2805_S), .p1(I_2869_D), .p2(I_3191_D));
	generic_cmos pass_157(.gn(I_93_S), .gp(I_95_D), .p1(I_575_S), .p2(I_319_D));
	generic_cmos pass_158(.gn(I_2807_S), .gp(I_2775_D), .p1(I_2871_D), .p2(I_2871_S));
	generic_cmos pass_159(.gn(I_2007_D), .gp(I_1973_D), .p1(I_2873_D), .p2(I_2969_D));
	generic_cmos pass_16(.gn(I_1099_S), .gp(I_1258_G), .p1(I_1227_D), .p2(I_1259_D));
	generic_cmos pass_160(.gn(I_395_D), .gp(I_329_D), .p1(I_293_D), .p2(I_293_S));
	generic_cmos pass_161(.gn(I_329_D), .gp(I_395_D), .p1(I_295_D), .p2(I_2329_D));
	generic_cmos pass_162(.gn(I_3265_S), .gp(I_3489_S), .p1(I_3169_S), .p2(I_3009_D));
	generic_cmos pass_163(.gn(I_2853_S), .gp(I_2791_S), .p1(I_2981_D), .p2(I_3013_D));
	generic_cmos pass_164(.gn(I_2791_S), .gp(I_2853_S), .p1(I_3013_S), .p2(I_3015_D));
	generic_cmos pass_165(.gn(I_3219_D), .gp(I_3059_D), .p1(I_3123_S), .p2(I_3027_D));
	generic_cmos pass_166(.gn(I_3191_S), .gp(I_3061_D), .p1(I_3125_S), .p2(I_3029_D));
	generic_cmos pass_167(.gn(I_3191_D), .gp(I_3063_D), .p1(I_3127_S), .p2(I_3031_D));
	generic_cmos pass_168(.gn(I_1973_D), .gp(I_2007_D), .p1(I_3993_S), .p2(I_3033_D));
	generic_cmos pass_169(.gn(I_3489_S), .gp(I_3265_S), .p1(I_3009_D), .p2(I_3073_D));
	generic_cmos pass_17(.gn(I_1045_D), .gp(I_789_D), .p1(I_2041_D), .p2(I_155_D));
	generic_cmos pass_170(.gn(I_2791_S), .gp(I_2853_S), .p1(I_3013_D), .p2(I_3013_S));
	generic_cmos pass_171(.gn(I_2853_S), .gp(I_2791_S), .p1(I_3015_D), .p2(I_3015_S));
	generic_cmos pass_172(.gn(I_3059_D), .gp(I_3219_D), .p1(I_3027_D), .p2(I_3985_D));
	generic_cmos pass_173(.gn(I_3061_D), .gp(I_3191_S), .p1(I_3029_D), .p2(I_3345_D));
	generic_cmos pass_174(.gn(I_3063_D), .gp(I_3191_D), .p1(I_3031_D), .p2(I_3031_S));
	generic_cmos pass_175(.gn(I_2007_D), .gp(I_1973_D), .p1(I_3033_D), .p2(I_3129_D));
	generic_cmos pass_176(.gn(I_251_S), .gp(I_315_D), .p1(I_311_D), .p2(I_375_D));
	generic_cmos pass_177(.gn(I_315_D), .gp(I_251_S), .p1(I_313_D), .p2(I_409_S));
	generic_cmos pass_178(.gn(I_3489_S), .gp(I_3265_S), .p1(I_3137_D), .p2(I_3169_D));
	generic_cmos pass_179(.gn(I_3013_S), .gp(I_2951_S), .p1(I_3141_D), .p2(I_3173_D));
	generic_cmos pass_18(.gn(I_1999_D), .gp(I_1297_D), .p1(I_1361_S), .p2(I_1265_D));
	generic_cmos pass_180(.gn(I_2951_S), .gp(I_3013_S), .p1(I_3173_S), .p2(I_3175_D));
	generic_cmos pass_181(.gn(I_3265_S), .gp(I_3489_S), .p1(I_3169_D), .p2(I_3169_S));
	generic_cmos pass_182(.gn(I_93_S), .gp(I_95_D), .p1(I_317_D), .p2(I_445_D));
	generic_cmos pass_183(.gn(I_2951_S), .gp(I_3013_S), .p1(I_3173_D), .p2(I_3173_S));
	generic_cmos pass_184(.gn(I_3013_S), .gp(I_2951_S), .p1(I_3175_D), .p2(I_3175_S));
	generic_cmos pass_185(.gn(I_3313_D), .gp(I_3345_S), .p1(I_3825_S), .p2(I_3185_S));
	generic_cmos pass_186(.gn(I_3985_D), .gp(I_3123_S), .p1(I_3219_D), .p2(I_3507_D));
	generic_cmos pass_187(.gn(I_3345_D), .gp(I_3125_S), .p1(I_3191_S), .p2(I_3189_S));
	generic_cmos pass_188(.gn(I_95_D), .gp(I_93_S), .p1(I_319_D), .p2(I_415_S));
	generic_cmos pass_189(.gn(I_3031_S), .gp(I_3127_S), .p1(I_3191_D), .p2(I_3191_S));
	generic_cmos pass_19(.gn(I_735_D), .gp(I_1301_D), .p1(I_1235_D), .p2(I_1267_D));
	generic_cmos pass_190(.gn(I_3555_G), .gp(I_3521_D), .p1(I_3489_S), .p2(I_3329_D));
	generic_cmos pass_191(.gn(I_3173_S), .gp(I_3111_S), .p1(I_3301_D), .p2(I_3333_D));
	generic_cmos pass_192(.gn(I_3111_S), .gp(I_3173_S), .p1(I_3333_S), .p2(I_3335_D));
	generic_cmos pass_193(.gn(I_3591_S), .gp(I_3369_D), .p1(I_3433_S), .p2(I_3337_D));
	generic_cmos pass_194(.gn(I_3499_D), .gp(I_3371_D), .p1(I_3435_S), .p2(I_3339_D));
	generic_cmos pass_195(.gn(I_3249_D), .gp(I_3281_S), .p1(I_3313_D), .p2(I_3345_D));
	generic_cmos pass_196(.gn(I_3507_D), .gp(I_3379_D), .p1(I_3443_S), .p2(I_3347_D));
	generic_cmos pass_197(.gn(I_3521_D), .gp(I_3555_G), .p1(I_3329_D), .p2(I_3393_D));
	generic_cmos pass_198(.gn(I_3111_S), .gp(I_3173_S), .p1(I_3333_D), .p2(I_3333_S));
	generic_cmos pass_199(.gn(I_3173_S), .gp(I_3111_S), .p1(I_3335_D), .p2(I_3335_S));
	generic_cmos pass_2(.gn(I_395_D), .gp(I_329_D), .p1(I_103_D), .p2(I_135_D));
	generic_cmos pass_20(.gn(I_1301_D), .gp(I_735_D), .p1(I_1237_D), .p2(I_1269_D));
	generic_cmos pass_200(.gn(I_3369_D), .gp(I_3591_S), .p1(I_3337_D), .p2(I_3499_D));
	generic_cmos pass_201(.gn(I_3371_D), .gp(I_3499_D), .p1(I_3339_D), .p2(I_3497_S));
	generic_cmos pass_202(.gn(I_3471_D), .gp(I_3503_S), .p1(I_3823_D), .p2(I_3535_D));
	generic_cmos pass_203(.gn(I_3281_S), .gp(I_3249_D), .p1(I_3345_D), .p2(I_3345_S));
	generic_cmos pass_204(.gn(I_3379_D), .gp(I_3507_D), .p1(I_3347_D), .p2(I_3503_D));
	generic_cmos pass_205(.gn(I_3521_D), .gp(I_3555_G), .p1(I_3457_D), .p2(I_3489_D));
	generic_cmos pass_206(.gn(I_3333_S), .gp(I_3271_S), .p1(I_3461_D), .p2(I_3493_D));
	generic_cmos pass_207(.gn(I_3271_S), .gp(I_3333_S), .p1(I_3493_S), .p2(I_3495_D));
	generic_cmos pass_208(.gn(I_3407_D), .gp(I_3439_S), .p1(I_3471_D), .p2(I_3503_D));
	generic_cmos pass_209(.gn(I_3555_G), .gp(I_3521_D), .p1(I_3489_D), .p2(I_3489_S));
	generic_cmos pass_21(.gn(I_315_D), .gp(I_251_S), .p1(I_1239_D), .p2(I_1271_D));
	generic_cmos pass_210(.gn(I_3271_S), .gp(I_3333_S), .p1(I_3493_D), .p2(I_3493_S));
	generic_cmos pass_211(.gn(I_3333_S), .gp(I_3271_S), .p1(I_3495_D), .p2(I_3495_S));
	generic_cmos pass_212(.gn(I_3499_D), .gp(I_3433_S), .p1(I_3591_S), .p2(I_3497_S));
	generic_cmos pass_213(.gn(I_3497_S), .gp(I_3435_S), .p1(I_3499_D), .p2(I_3499_S));
	generic_cmos pass_214(.gn(I_3439_S), .gp(I_3407_D), .p1(I_3503_D), .p2(I_3503_S));
	generic_cmos pass_215(.gn(I_3503_D), .gp(I_3443_S), .p1(I_3507_D), .p2(I_3827_D));
	generic_cmos pass_216(.gn(I_3493_S), .gp(I_3431_S), .p1(I_3621_D), .p2(I_3653_D));
	generic_cmos pass_217(.gn(I_3431_S), .gp(I_3493_S), .p1(I_3653_S), .p2(I_3655_D));
	generic_cmos pass_218(.gn(I_3823_D), .gp(I_3695_D), .p1(I_3759_S), .p2(I_3663_D));
	generic_cmos pass_219(.gn(I_3827_D), .gp(I_3699_D), .p1(I_3763_S), .p2(I_3667_D));
	generic_cmos pass_22(.gn(I_1469_D), .gp(I_1213_D), .p1(I_1247_D), .p2(I_1279_D));
	generic_cmos pass_220(.gn(I_3829_D), .gp(I_3701_D), .p1(I_3765_S), .p2(I_3669_D));
	generic_cmos pass_221(.gn(I_3431_S), .gp(I_3493_S), .p1(I_3653_D), .p2(I_3653_S));
	generic_cmos pass_222(.gn(I_3493_S), .gp(I_3431_S), .p1(I_3655_D), .p2(I_3655_S));
	generic_cmos pass_223(.gn(I_3695_D), .gp(I_3823_D), .p1(I_3663_D), .p2(I_3663_S));
	generic_cmos pass_224(.gn(I_3699_D), .gp(I_3827_D), .p1(I_3667_D), .p2(I_3667_S));
	generic_cmos pass_225(.gn(I_3701_D), .gp(I_3829_D), .p1(I_3669_D), .p2(I_3669_S));
	generic_cmos pass_226(.gn(I_3653_S), .gp(I_3591_S), .p1(I_3781_D), .p2(I_3813_D));
	generic_cmos pass_227(.gn(I_3591_S), .gp(I_3653_S), .p1(I_3813_S), .p2(I_3815_D));
	generic_cmos pass_228(.gn(I_3591_S), .gp(I_3653_S), .p1(I_3813_D), .p2(I_3813_S));
	generic_cmos pass_229(.gn(I_3653_S), .gp(I_3591_S), .p1(I_3815_D), .p2(I_3815_S));
	generic_cmos pass_23(.gn(I_93_S), .gp(I_95_D), .p1(I_477_D), .p2(I_157_D));
	generic_cmos pass_230(.gn(I_3663_S), .gp(I_3759_S), .p1(I_3823_D), .p2(I_3823_S));
	generic_cmos pass_231(.gn(I_3953_D), .gp(I_3985_S), .p1(I_3825_D), .p2(I_3825_S));
	generic_cmos pass_232(.gn(I_3667_S), .gp(I_3763_S), .p1(I_3827_D), .p2(I_3829_D));
	generic_cmos pass_233(.gn(I_3669_S), .gp(I_3765_S), .p1(I_3829_D), .p2(I_3829_S));
	generic_cmos pass_234(.gn(I_3889_D), .gp(I_3921_S), .p1(I_3953_D), .p2(I_3985_D));
	generic_cmos pass_235(.gn(I_3921_S), .gp(I_3889_D), .p1(I_3985_D), .p2(I_3985_S));
	generic_cmos pass_236(.gn(I_329_D), .gp(I_395_D), .p1(I_421_D), .p2(I_453_D));
	generic_cmos pass_237(.gn(I_395_D), .gp(I_329_D), .p1(I_423_D), .p2(I_455_D));
	generic_cmos pass_238(.gn(I_251_S), .gp(I_315_D), .p1(I_439_D), .p2(I_471_D));
	generic_cmos pass_239(.gn(I_315_D), .gp(I_251_S), .p1(I_475_D), .p2(I_473_D));
	generic_cmos pass_24(.gn(I_715_D), .gp(I_1097_S), .p1(I_1253_D), .p2(I_1253_S));
	generic_cmos pass_240(.gn(I_789_D), .gp(I_1045_D), .p1(I_443_D), .p2(I_475_D));
	generic_cmos pass_241(.gn(I_509_D), .gp(I_573_D), .p1(I_445_D), .p2(I_477_D));
	generic_cmos pass_242(.gn(I_95_D), .gp(I_93_S), .p1(I_447_D), .p2(I_479_D));
	generic_cmos pass_243(.gn(I_395_D), .gp(I_329_D), .p1(I_453_D), .p2(I_453_S));
	generic_cmos pass_244(.gn(I_329_D), .gp(I_395_D), .p1(I_455_D), .p2(I_1415_S));
	generic_cmos pass_245(.gn(I_315_D), .gp(I_251_S), .p1(I_471_D), .p2(I_471_S));
	generic_cmos pass_246(.gn(I_251_S), .gp(I_315_D), .p1(I_473_D), .p2(I_505_D));
	generic_cmos pass_247(.gn(I_1045_D), .gp(I_789_D), .p1(I_475_D), .p2(I_2201_D));
	generic_cmos pass_248(.gn(I_573_D), .gp(I_509_D), .p1(I_477_D), .p2(I_477_S));
	generic_cmos pass_249(.gn(I_93_S), .gp(I_95_D), .p1(I_479_D), .p2(I_575_S));
	generic_cmos pass_25(.gn(I_1097_S), .gp(I_715_D), .p1(I_1255_D), .p2(I_2329_D));
	generic_cmos pass_250(.gn(I_393_S), .gp(I_555_D), .p1(I_581_D), .p2(I_613_D));
	generic_cmos pass_251(.gn(I_555_D), .gp(I_393_S), .p1(I_583_D), .p2(I_615_D));
	generic_cmos pass_252(.gn(I_1045_D), .gp(I_789_D), .p1(I_2841_D), .p2(I_631_D));
	generic_cmos pass_253(.gn(I_251_S), .gp(I_315_D), .p1(I_601_D), .p2(I_633_D));
	generic_cmos pass_254(.gn(I_93_S), .gp(I_95_D), .p1(I_957_D), .p2(I_637_D));
	generic_cmos pass_255(.gn(I_555_D), .gp(I_393_S), .p1(I_613_D), .p2(I_613_S));
	generic_cmos pass_256(.gn(I_393_S), .gp(I_555_D), .p1(I_615_D), .p2(I_2169_D));
	generic_cmos pass_257(.gn(I_789_D), .gp(I_1045_D), .p1(I_631_D), .p2(I_727_D));
	generic_cmos pass_258(.gn(I_315_D), .gp(I_251_S), .p1(I_633_D), .p2(I_729_S));
	generic_cmos pass_259(.gn(I_95_D), .gp(I_93_S), .p1(I_637_D), .p2(I_733_S));
	generic_cmos pass_26(.gn(I_1099_S), .gp(I_1258_G), .p1(I_1257_D), .p2(I_1355_D));
	generic_cmos pass_260(.gn(I_93_S), .gp(I_95_D), .p1(I_1407_D), .p2(I_639_S));
	generic_cmos pass_261(.gn(I_393_S), .gp(I_555_D), .p1(I_741_D), .p2(I_773_D));
	generic_cmos pass_262(.gn(I_555_D), .gp(I_393_S), .p1(I_743_D), .p2(I_775_D));
	generic_cmos pass_263(.gn(I_713_S), .gp(I_779_S), .p1(I_1415_S), .p2(I_777_D));
	generic_cmos pass_264(.gn(I_315_D), .gp(I_251_S), .p1(I_759_D), .p2(I_791_D));
	generic_cmos pass_265(.gn(I_315_D), .gp(I_251_S), .p1(I_795_D), .p2(I_793_D));
	generic_cmos pass_266(.gn(I_789_D), .gp(I_1045_D), .p1(I_763_D), .p2(I_795_D));
	generic_cmos pass_267(.gn(I_95_D), .gp(I_93_S), .p1(I_765_D), .p2(I_797_D));
	generic_cmos pass_268(.gn(I_555_D), .gp(I_393_S), .p1(I_773_D), .p2(I_773_S));
	generic_cmos pass_269(.gn(I_393_S), .gp(I_555_D), .p1(I_775_D), .p2(I_2329_D));
	generic_cmos pass_27(.gn(I_1258_G), .gp(I_1099_S), .p1(I_1259_D), .p2(I_1259_S));
	generic_cmos pass_270(.gn(I_779_S), .gp(I_713_S), .p1(I_777_D), .p2(I_873_D));
	generic_cmos pass_271(.gn(I_251_S), .gp(I_315_D), .p1(I_791_D), .p2(I_855_D));
	generic_cmos pass_272(.gn(I_251_S), .gp(I_315_D), .p1(I_793_D), .p2(I_825_D));
	generic_cmos pass_273(.gn(I_1045_D), .gp(I_789_D), .p1(I_795_D), .p2(I_2361_D));
	generic_cmos pass_274(.gn(I_93_S), .gp(I_95_D), .p1(I_797_D), .p2(I_925_D));
	generic_cmos pass_275(.gn(I_93_S), .gp(I_95_D), .p1(I_1407_D), .p2(I_799_S));
	generic_cmos pass_276(.gn(I_393_S), .gp(I_555_D), .p1(I_901_D), .p2(I_933_D));
	generic_cmos pass_277(.gn(I_555_D), .gp(I_393_S), .p1(I_903_D), .p2(I_935_D));
	generic_cmos pass_278(.gn(I_713_S), .gp(I_779_S), .p1(I_2329_D), .p2(I_937_D));
	generic_cmos pass_279(.gn(I_251_S), .gp(I_315_D), .p1(I_919_D), .p2(I_951_D));
	generic_cmos pass_28(.gn(I_1297_D), .gp(I_1999_D), .p1(I_1265_D), .p2(I_2071_S));
	generic_cmos pass_280(.gn(I_251_S), .gp(I_315_D), .p1(I_921_D), .p2(I_953_D));
	generic_cmos pass_281(.gn(I_735_D), .gp(I_989_D), .p1(I_925_D), .p2(I_957_D));
	generic_cmos pass_282(.gn(I_93_S), .gp(I_95_D), .p1(I_1279_D), .p2(I_959_D));
	generic_cmos pass_283(.gn(I_555_D), .gp(I_393_S), .p1(I_933_D), .p2(I_933_S));
	generic_cmos pass_284(.gn(I_393_S), .gp(I_555_D), .p1(I_935_D), .p2(I_1415_S));
	generic_cmos pass_285(.gn(I_779_S), .gp(I_713_S), .p1(I_937_D), .p2(I_1033_D));
	generic_cmos pass_286(.gn(I_315_D), .gp(I_251_S), .p1(I_951_D), .p2(I_1111_D));
	generic_cmos pass_287(.gn(I_315_D), .gp(I_251_S), .p1(I_953_D), .p2(I_1049_S));
	generic_cmos pass_288(.gn(I_989_D), .gp(I_735_D), .p1(I_957_D), .p2(I_957_S));
	generic_cmos pass_289(.gn(I_95_D), .gp(I_93_S), .p1(I_959_D), .p2(I_1055_S));
	generic_cmos pass_29(.gn(I_1301_D), .gp(I_735_D), .p1(I_1267_D), .p2(I_1267_S));
	generic_cmos pass_3(.gn(I_1097_S), .gp(I_715_D), .p1(I_1061_D), .p2(I_1093_D));
	generic_cmos pass_30(.gn(I_735_D), .gp(I_1301_D), .p1(I_1269_D), .p2(I_1269_S));
	generic_cmos pass_31(.gn(I_251_S), .gp(I_315_D), .p1(I_1271_D), .p2(I_1335_D));
	generic_cmos pass_32(.gn(I_1213_D), .gp(I_1469_D), .p1(I_1279_D), .p2(I_1279_S));
	generic_cmos pass_33(.gn(I_395_D), .gp(I_329_D), .p1(I_133_D), .p2(I_133_S));
	generic_cmos pass_34(.gn(I_329_D), .gp(I_395_D), .p1(I_135_D), .p2(I_2169_D));
	generic_cmos pass_35(.gn(I_1097_S), .gp(I_715_D), .p1(I_1381_D), .p2(I_1413_D));
	generic_cmos pass_36(.gn(I_715_D), .gp(I_1097_S), .p1(I_1383_D), .p2(I_1415_D));
	generic_cmos pass_37(.gn(I_1101_S), .gp(I_1420_S), .p1(I_1385_D), .p2(I_1417_D));
	generic_cmos pass_38(.gn(I_1420_S), .gp(I_1101_S), .p1(I_1387_D), .p2(I_1419_D));
	generic_cmos pass_39(.gn(I_1589_S), .gp(I_1749_S), .p1(I_1525_D), .p2(I_1427_D));
	generic_cmos pass_4(.gn(I_715_D), .gp(I_1097_S), .p1(I_1063_D), .p2(I_1095_D));
	generic_cmos pass_40(.gn(I_1749_S), .gp(I_1589_S), .p1(I_1397_D), .p2(I_1429_D));
	generic_cmos pass_41(.gn(I_251_S), .gp(I_315_D), .p1(I_1399_D), .p2(I_1431_D));
	generic_cmos pass_42(.gn(I_789_D), .gp(I_1045_D), .p1(I_1401_D), .p2(I_1433_D));
	generic_cmos pass_43(.gn(I_93_S), .gp(I_95_D), .p1(I_1407_D), .p2(I_1439_D));
	generic_cmos pass_44(.gn(I_715_D), .gp(I_1097_S), .p1(I_1413_D), .p2(I_1413_S));
	generic_cmos pass_45(.gn(I_1097_S), .gp(I_715_D), .p1(I_1415_D), .p2(I_1415_S));
	generic_cmos pass_46(.gn(I_1420_S), .gp(I_1101_S), .p1(I_1417_D), .p2(I_1417_S));
	generic_cmos pass_47(.gn(I_1101_S), .gp(I_1420_S), .p1(I_1419_D), .p2(I_1419_S));
	generic_cmos pass_48(.gn(I_2071_S), .gp(I_1361_S), .p1(I_1999_D), .p2(I_1425_S));
	generic_cmos pass_49(.gn(I_1749_S), .gp(I_1589_S), .p1(I_1427_D), .p2(I_1523_S));
	generic_cmos pass_5(.gn(I_1045_D), .gp(I_789_D), .p1(I_2681_D), .p2(I_1111_D));
	generic_cmos pass_50(.gn(I_1589_S), .gp(I_1749_S), .p1(I_1429_D), .p2(I_1461_D));
	generic_cmos pass_51(.gn(I_315_D), .gp(I_251_S), .p1(I_1431_D), .p2(I_1433_D));
	generic_cmos pass_52(.gn(I_1045_D), .gp(I_789_D), .p1(I_1433_D), .p2(I_2521_D));
	generic_cmos pass_53(.gn(I_95_D), .gp(I_93_S), .p1(I_1439_D), .p2(I_1439_S));
	generic_cmos pass_54(.gn(I_251_S), .gp(I_315_D), .p1(I_153_D), .p2(I_185_D));
	generic_cmos pass_55(.gn(I_1671_S), .gp(I_1411_S), .p1(I_1537_D), .p2(I_1569_D));
	generic_cmos pass_56(.gn(I_1411_S), .gp(I_1671_S), .p1(I_1539_D), .p2(I_1571_D));
	generic_cmos pass_57(.gn(I_1576_S), .gp(I_1051_S), .p1(I_1541_D), .p2(I_1573_D));
	generic_cmos pass_58(.gn(I_1051_S), .gp(I_1576_S), .p1(I_1573_S), .p2(I_1575_D));
	generic_cmos pass_59(.gn(I_789_D), .gp(I_1045_D), .p1(I_155_D), .p2(VSS));
	generic_cmos pass_6(.gn(I_95_D), .gp(I_93_S), .p1(I_1087_D), .p2(I_1119_D));
	generic_cmos pass_60(.gn(I_1623_D), .gp(I_1753_S), .p1(I_1559_D), .p2(I_1591_D));
	generic_cmos pass_61(.gn(I_1753_S), .gp(I_1623_D), .p1(I_1561_D), .p2(I_1593_D));
	generic_cmos pass_62(.gn(I_1411_S), .gp(I_1671_S), .p1(I_1569_D), .p2(I_1891_S));
	generic_cmos pass_63(.gn(I_95_D), .gp(I_93_S), .p1(I_157_D), .p2(I_253_S));
	generic_cmos pass_64(.gn(I_1671_S), .gp(I_1411_S), .p1(I_1571_D), .p2(I_1571_S));
	generic_cmos pass_65(.gn(I_1051_S), .gp(I_1576_S), .p1(I_1573_D), .p2(I_1573_S));
	generic_cmos pass_66(.gn(I_1576_S), .gp(I_1051_S), .p1(I_1575_D), .p2(I_1575_S));
	generic_cmos pass_67(.gn(I_93_S), .gp(I_95_D), .p1(I_1407_D), .p2(I_159_S));
	generic_cmos pass_68(.gn(I_1753_S), .gp(I_1623_D), .p1(I_1591_D), .p2(I_1845_D));
	generic_cmos pass_69(.gn(I_1623_D), .gp(I_1753_S), .p1(I_1593_D), .p2(I_1593_S));
	generic_cmos pass_7(.gn(I_715_D), .gp(I_1097_S), .p1(I_1093_D), .p2(I_1093_S));
	generic_cmos pass_70(.gn(I_1730_G), .gp(I_1761_D), .p1(I_1697_D), .p2(I_1729_D));
	generic_cmos pass_71(.gn(I_1761_D), .gp(I_1730_G), .p1(I_1699_D), .p2(I_1731_D));
	generic_cmos pass_72(.gn(I_1573_S), .gp(I_1511_S), .p1(I_1701_D), .p2(I_1733_D));
	generic_cmos pass_73(.gn(I_1511_S), .gp(I_1573_S), .p1(I_1733_S), .p2(I_1735_D));
	generic_cmos pass_74(.gn(I_1761_D), .gp(I_1730_G), .p1(I_1729_D), .p2(I_1729_S));
	generic_cmos pass_75(.gn(I_1730_G), .gp(I_1761_D), .p1(I_1731_D), .p2(I_1731_S));
	generic_cmos pass_76(.gn(I_1511_S), .gp(I_1573_S), .p1(I_1733_D), .p2(I_1733_S));
	generic_cmos pass_77(.gn(I_1573_S), .gp(I_1511_S), .p1(I_1735_D), .p2(I_1735_S));
	generic_cmos pass_78(.gn(I_1733_S), .gp(I_1671_S), .p1(I_1861_D), .p2(I_1893_D));
	generic_cmos pass_79(.gn(I_1671_S), .gp(I_1733_S), .p1(I_1893_S), .p2(I_1895_D));
	generic_cmos pass_8(.gn(I_1097_S), .gp(I_715_D), .p1(I_1095_D), .p2(I_2169_D));
	generic_cmos pass_80(.gn(I_1908_S), .gp(I_503_D), .p1(I_1879_D), .p2(I_1911_D));
	generic_cmos pass_81(.gn(I_503_D), .gp(I_1908_S), .p1(I_1881_D), .p2(I_1913_D));
	generic_cmos pass_82(.gn(I_1671_S), .gp(I_1733_S), .p1(I_1893_D), .p2(I_1893_S));
	generic_cmos pass_83(.gn(I_1733_S), .gp(I_1671_S), .p1(I_1895_D), .p2(I_1895_S));
	generic_cmos pass_84(.gn(I_2033_D), .gp(I_2065_S), .p1(I_2545_S), .p2(I_1906_S));
	generic_cmos pass_85(.gn(I_503_D), .gp(I_1908_S), .p1(I_1911_D), .p2(I_1911_S));
	generic_cmos pass_86(.gn(I_1908_S), .gp(I_503_D), .p1(I_1913_D), .p2(I_1913_S));
	generic_cmos pass_87(.gn(I_2305_S), .gp(I_2529_S), .p1(I_2209_S), .p2(I_2049_D));
	generic_cmos pass_88(.gn(I_1893_S), .gp(I_1831_S), .p1(I_2021_D), .p2(I_2053_D));
	generic_cmos pass_89(.gn(I_1831_S), .gp(I_1893_S), .p1(I_2053_S), .p2(I_2055_D));
	generic_cmos pass_9(.gn(I_789_D), .gp(I_1045_D), .p1(I_1111_D), .p2(I_1207_D));
	generic_cmos pass_90(.gn(I_1969_D), .gp(I_2001_S), .p1(I_2033_D), .p2(I_2709_S));
	generic_cmos pass_91(.gn(I_2231_D), .gp(I_2103_D), .p1(I_2167_S), .p2(I_2071_D));
	generic_cmos pass_92(.gn(I_1973_D), .gp(I_2007_D), .p1(I_2041_D), .p2(I_2073_D));
	generic_cmos pass_93(.gn(I_2529_S), .gp(I_2305_S), .p1(I_2049_D), .p2(I_2113_D));
	generic_cmos pass_94(.gn(I_1831_S), .gp(I_1893_S), .p1(I_2053_D), .p2(I_2053_S));
	generic_cmos pass_95(.gn(I_1893_S), .gp(I_1831_S), .p1(I_2055_D), .p2(I_2055_S));
	generic_cmos pass_96(.gn(I_2001_S), .gp(I_1969_D), .p1(I_2709_S), .p2(I_2065_S));
	generic_cmos pass_97(.gn(I_2103_D), .gp(I_2231_D), .p1(I_2071_D), .p2(I_2071_S));
	generic_cmos pass_98(.gn(I_2007_D), .gp(I_1973_D), .p1(I_2073_D), .p2(I_2169_D));
	generic_cmos pass_99(.gn(I_2529_S), .gp(I_2305_S), .p1(I_2177_D), .p2(I_2209_D));

endmodule

